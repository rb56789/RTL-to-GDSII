`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:PhD 
// Engineer:ANURAJ V 
// 
// Create Date: 03/20/2024 09:35:02 PM
// Design Name: 
// Module Name: WA_32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module FA(a,b,cin,sum,carry);
    input a,b,cin;
    output sum,carry;
    
wire [2:0] faw;     

xor(faw[0],a,b);
xor(sum,faw[0],cin);        

and(faw[1],a,b);
and(faw[2],faw[0],cin);

or(carry,faw[1],faw[2]);    
endmodule

module HA(a,b,sum_h,carry_h);
    input a,b;
    output sum_h,carry_h;
 xor(sum_h, a, b);
 and(carry_h, a, b);
endmodule

module WA_32(x,y,z);
input [31:0] x,y;
output [64:0] z;

//wire [62:0] p;
wire [160:0] hca;
wire [160:0] hsu;
wire [960:0] fca;
wire [960:0] fsu;

    reg[31:0] pp[31:0];
    integer i, j;

    always @(x, y) begin
        for(i = 0;i < 32;i = i+1)
            for(j = 0;j < 32;j = j+1)
                pp[i][j] = x[i] & y[j];
    end

assign z[0] = pp[0][0];

//1st stage
HA HA1 (.a(pp[1][0]),.b(pp[0][1]),.sum_h(z[1]),.carry_h(hca[1]));//p1
FA FA1 (.a(pp[2][0]),.b(pp[1][1]),.cin(pp[0][2]),.sum(fsu[1]),.carry(fca[1]));
FA FA2 (.a(pp[3][0]),.b(pp[2][1]),.cin(pp[1][2]),.sum(fsu[2]),.carry(fca[2]));
FA FA3 (.a(pp[4][0]),.b(pp[3][1]),.cin(pp[2][2]),.sum(fsu[3]),.carry(fca[3]));
HA HA2 (.a(pp[1][3]),.b(pp[0][4]),.sum_h(hsu[2]),.carry_h(hca[2]));
FA FA4 (.a(pp[5][0]),.b(pp[4][1]),.cin(pp[3][2]),.sum(fsu[4]),.carry(fca[4]));
FA FA5 (.a(pp[2][3]),.b(pp[1][4]),.cin(pp[0][5]),.sum(fsu[5]),.carry(fca[5]));
FA FA6 (.a(pp[6][0]),.b(pp[5][1]),.cin(pp[4][2]),.sum(fsu[6]),.carry(fca[6]));
FA FA7 (.a(pp[3][3]),.b(pp[2][4]),.cin(pp[1][5]),.sum(fsu[7]),.carry(fca[7]));
FA FA8 (.a(pp[7][0]),.b(pp[6][1]),.cin(pp[5][2]),.sum(fsu[8]),.carry(fca[8]));
FA FA9 (.a(pp[4][3]),.b(pp[3][4]),.cin(pp[2][5]),.sum(fsu[9]),.carry(fca[9]));
HA HA3 (.a(pp[1][6]),.b(pp[0][7]),.sum_h(hsu[3]),.carry_h(hca[3]));
FA FA10 (.a(pp[8][0]),.b(pp[7][1]),.cin(pp[6][2]),.sum(fsu[10]),.carry(fca[10]));
FA FA11 (.a(pp[5][3]),.b(pp[4][4]),.cin(pp[3][5]),.sum(fsu[11]),.carry(fca[11]));
FA FA12 (.a(pp[2][6]),.b(pp[1][7]),.cin(pp[0][8]),.sum(fsu[12]),.carry(fca[12]));
FA FA13 (.a(pp[9][0]),.b(pp[8][1]),.cin(pp[7][2]),.sum(fsu[13]),.carry(fca[13]));
FA FA14 (.a(pp[6][3]),.b(pp[5][4]),.cin(pp[4][5]),.sum(fsu[14]),.carry(fca[14]));
FA FA15 (.a(pp[3][6]),.b(pp[2][7]),.cin(pp[1][8]),.sum(fsu[15]),.carry(fca[15]));
FA FA16 (.a(pp[10][0]),.b(pp[9][1]),.cin(pp[8][2]),.sum(fsu[16]),.carry(fca[16]));
FA FA17 (.a(pp[7][3]),.b(pp[6][4]),.cin(pp[5][5]),.sum(fsu[17]),.carry(fca[17]));
FA FA18 (.a(pp[4][6]),.b(pp[3][7]),.cin(pp[2][8]),.sum(fsu[18]),.carry(fca[18]));
HA HA4 (.a(pp[1][9]),.b(pp[0][10]),.sum_h(hsu[4]),.carry_h(hca[4]));
FA FA19 (.a(pp[11][0]),.b(pp[10][1]),.cin(pp[9][2]),.sum(fsu[19]),.carry(fca[19]));
FA FA20 (.a(pp[8][3]),.b(pp[7][4]),.cin(pp[6][5]),.sum(fsu[20]),.carry(fca[20]));
FA FA21 (.a(pp[5][6]),.b(pp[4][7]),.cin(pp[3][8]),.sum(fsu[21]),.carry(fca[21]));
FA FA22 (.a(pp[2][9]),.b(pp[1][10]),.cin(pp[0][11]),.sum(fsu[22]),.carry(fca[22]));
FA FA23 (.a(pp[12][0]),.b(pp[11][1]),.cin(pp[10][2]),.sum(fsu[23]),.carry(fca[23]));
FA FA24 (.a(pp[9][3]),.b(pp[8][4]),.cin(pp[7][5]),.sum(fsu[24]),.carry(fca[24]));
FA FA25 (.a(pp[6][6]),.b(pp[5][7]),.cin(pp[4][8]),.sum(fsu[25]),.carry(fca[25]));
FA FA26 (.a(pp[3][9]),.b(pp[2][10]),.cin(pp[1][11]),.sum(fsu[26]),.carry(fca[26]));
FA FA27 (.a(pp[13][0]),.b(pp[12][1]),.cin(pp[11][2]),.sum(fsu[27]),.carry(fca[27]));
FA FA28 (.a(pp[10][3]),.b(pp[9][4]),.cin(pp[8][5]),.sum(fsu[28]),.carry(fca[28]));
FA FA29 (.a(pp[7][6]),.b(pp[6][7]),.cin(pp[5][8]),.sum(fsu[29]),.carry(fca[29]));
FA FA30 (.a(pp[4][9]),.b(pp[3][10]),.cin(pp[2][11]),.sum(fsu[30]),.carry(fca[30]));
HA HA5 (.a(pp[1][12]),.b(pp[0][13]),.sum_h(hsu[5]),.carry_h(hca[5]));
FA FA31 (.a(pp[14][0]),.b(pp[13][1]),.cin(pp[12][2]),.sum(fsu[31]),.carry(fca[31]));
FA FA32 (.a(pp[11][3]),.b(pp[10][4]),.cin(pp[9][5]),.sum(fsu[32]),.carry(fca[32]));
FA FA33 (.a(pp[8][6]),.b(pp[7][7]),.cin(pp[6][8]),.sum(fsu[33]),.carry(fca[33]));
FA FA34 (.a(pp[5][9]),.b(pp[4][10]),.cin(pp[3][11]),.sum(fsu[34]),.carry(fca[34]));
FA FA35 (.a(pp[2][12]),.b(pp[1][13]),.cin(pp[0][14]),.sum(fsu[35]),.carry(fca[35]));
FA FA36 (.a(pp[15][0]),.b(pp[14][1]),.cin(pp[13][2]),.sum(fsu[36]),.carry(fca[36]));
FA FA37 (.a(pp[12][3]),.b(pp[11][4]),.cin(pp[10][5]),.sum(fsu[37]),.carry(fca[37]));
FA FA38 (.a(pp[9][6]),.b(pp[8][7]),.cin(pp[7][8]),.sum(fsu[38]),.carry(fca[38]));
FA FA39 (.a(pp[6][9]),.b(pp[5][10]),.cin(pp[4][11]),.sum(fsu[39]),.carry(fca[39]));
FA FA40 (.a(pp[3][12]),.b(pp[2][13]),.cin(pp[1][14]),.sum(fsu[40]),.carry(fca[40]));
FA FA41 (.a(pp[16][0]),.b(pp[15][1]),.cin(pp[14][2]),.sum(fsu[41]),.carry(fca[41]));
FA FA42 (.a(pp[13][3]),.b(pp[12][4]),.cin(pp[11][5]),.sum(fsu[42]),.carry(fca[42]));
FA FA43 (.a(pp[10][6]),.b(pp[9][7]),.cin(pp[8][8]),.sum(fsu[43]),.carry(fca[43]));
FA FA44 (.a(pp[7][9]),.b(pp[6][10]),.cin(pp[5][11]),.sum(fsu[44]),.carry(fca[44]));
FA FA45 (.a(pp[4][12]),.b(pp[3][13]),.cin(pp[2][14]),.sum(fsu[45]),.carry(fca[45]));
HA HA6 (.a(pp[1][15]),.b(pp[0][16]),.sum_h(hsu[6]),.carry_h(hca[6]));
FA FA46 (.a(pp[17][0]),.b(pp[16][1]),.cin(pp[15][2]),.sum(fsu[46]),.carry(fca[46]));
FA FA47 (.a(pp[14][3]),.b(pp[13][4]),.cin(pp[12][5]),.sum(fsu[47]),.carry(fca[47]));
FA FA48 (.a(pp[11][6]),.b(pp[10][7]),.cin(pp[9][8]),.sum(fsu[48]),.carry(fca[48]));
FA FA49 (.a(pp[8][9]),.b(pp[7][10]),.cin(pp[6][11]),.sum(fsu[49]),.carry(fca[49]));
FA FA50 (.a(pp[5][12]),.b(pp[4][13]),.cin(pp[3][14]),.sum(fsu[50]),.carry(fca[50]));
FA FA51 (.a(pp[2][15]),.b(pp[1][16]),.cin(pp[0][17]),.sum(fsu[51]),.carry(fca[51]));
FA FA52 (.a(pp[18][0]),.b(pp[17][1]),.cin(pp[16][2]),.sum(fsu[52]),.carry(fca[52]));
FA FA53 (.a(pp[15][3]),.b(pp[14][4]),.cin(pp[13][5]),.sum(fsu[53]),.carry(fca[53]));
FA FA54 (.a(pp[12][6]),.b(pp[11][7]),.cin(pp[10][8]),.sum(fsu[54]),.carry(fca[54]));
FA FA55 (.a(pp[9][9]),.b(pp[8][10]),.cin(pp[7][11]),.sum(fsu[55]),.carry(fca[55]));
FA FA56 (.a(pp[6][12]),.b(pp[5][13]),.cin(pp[4][14]),.sum(fsu[56]),.carry(fca[56]));
FA FA57 (.a(pp[3][15]),.b(pp[2][16]),.cin(pp[1][17]),.sum(fsu[57]),.carry(fca[57]));
FA FA58 (.a(pp[19][0]),.b(pp[18][1]),.cin(pp[17][2]),.sum(fsu[58]),.carry(fca[58]));
FA FA59 (.a(pp[16][3]),.b(pp[15][4]),.cin(pp[14][5]),.sum(fsu[59]),.carry(fca[59]));
FA FA60 (.a(pp[13][6]),.b(pp[12][7]),.cin(pp[11][8]),.sum(fsu[60]),.carry(fca[60]));
FA FA61 (.a(pp[10][9]),.b(pp[9][10]),.cin(pp[8][11]),.sum(fsu[61]),.carry(fca[61]));
FA FA62 (.a(pp[7][12]),.b(pp[6][13]),.cin(pp[5][14]),.sum(fsu[62]),.carry(fca[62]));
FA FA63 (.a(pp[4][15]),.b(pp[3][16]),.cin(pp[2][17]),.sum(fsu[63]),.carry(fca[63]));
HA HA7 (.a(pp[1][18]),.b(pp[0][19]),.sum_h(hsu[7]),.carry_h(hca[7]));
FA FA64 (.a(pp[20][0]),.b(pp[19][1]),.cin(pp[18][2]),.sum(fsu[64]),.carry(fca[64]));
FA FA65 (.a(pp[17][3]),.b(pp[16][4]),.cin(pp[15][5]),.sum(fsu[65]),.carry(fca[65]));
FA FA66 (.a(pp[14][6]),.b(pp[13][7]),.cin(pp[12][8]),.sum(fsu[66]),.carry(fca[66]));
FA FA67 (.a(pp[11][9]),.b(pp[10][10]),.cin(pp[9][11]),.sum(fsu[67]),.carry(fca[67]));
FA FA68 (.a(pp[8][12]),.b(pp[7][13]),.cin(pp[6][14]),.sum(fsu[68]),.carry(fca[68]));
FA FA69 (.a(pp[5][15]),.b(pp[4][16]),.cin(pp[3][17]),.sum(fsu[69]),.carry(fca[69]));
FA FA70 (.a(pp[2][18]),.b(pp[1][19]),.cin(pp[0][20]),.sum(fsu[70]),.carry(fca[70]));
FA FA71 (.a(pp[21][0]),.b(pp[20][1]),.cin(pp[19][2]),.sum(fsu[71]),.carry(fca[71]));
FA FA72 (.a(pp[18][3]),.b(pp[17][4]),.cin(pp[16][5]),.sum(fsu[72]),.carry(fca[72]));
FA FA73 (.a(pp[15][6]),.b(pp[14][7]),.cin(pp[13][8]),.sum(fsu[73]),.carry(fca[73]));
FA FA74 (.a(pp[12][9]),.b(pp[11][10]),.cin(pp[10][11]),.sum(fsu[74]),.carry(fca[74]));
FA FA75 (.a(pp[9][12]),.b(pp[8][13]),.cin(pp[7][14]),.sum(fsu[75]),.carry(fca[75]));
FA FA76 (.a(pp[6][15]),.b(pp[5][16]),.cin(pp[4][17]),.sum(fsu[76]),.carry(fca[76]));
FA FA77 (.a(pp[3][18]),.b(pp[2][19]),.cin(pp[1][20]),.sum(fsu[77]),.carry(fca[77]));
FA FA78 (.a(pp[22][0]),.b(pp[21][1]),.cin(pp[20][2]),.sum(fsu[78]),.carry(fca[78]));
FA FA79 (.a(pp[19][3]),.b(pp[18][4]),.cin(pp[17][5]),.sum(fsu[79]),.carry(fca[79]));
FA FA80 (.a(pp[16][6]),.b(pp[15][7]),.cin(pp[14][8]),.sum(fsu[80]),.carry(fca[80]));
FA FA81 (.a(pp[13][9]),.b(pp[12][10]),.cin(pp[11][11]),.sum(fsu[81]),.carry(fca[81]));
FA FA82 (.a(pp[10][12]),.b(pp[9][13]),.cin(pp[8][14]),.sum(fsu[82]),.carry(fca[82]));
FA FA83 (.a(pp[7][15]),.b(pp[6][16]),.cin(pp[5][17]),.sum(fsu[83]),.carry(fca[83]));
FA FA84 (.a(pp[4][18]),.b(pp[3][19]),.cin(pp[2][20]),.sum(fsu[84]),.carry(fca[84]));
HA HA8 (.a(pp[1][21]),.b(pp[0][22]),.sum_h(hsu[8]),.carry_h(hca[8]));
FA FA85 (.a(pp[23][0]),.b(pp[22][1]),.cin(pp[21][2]),.sum(fsu[85]),.carry(fca[85]));
FA FA86 (.a(pp[20][3]),.b(pp[19][4]),.cin(pp[18][5]),.sum(fsu[86]),.carry(fca[86]));
FA FA87 (.a(pp[17][6]),.b(pp[16][7]),.cin(pp[15][8]),.sum(fsu[87]),.carry(fca[87]));
FA FA88 (.a(pp[14][9]),.b(pp[13][10]),.cin(pp[12][11]),.sum(fsu[88]),.carry(fca[88]));
FA FA89 (.a(pp[11][12]),.b(pp[10][13]),.cin(pp[9][14]),.sum(fsu[89]),.carry(fca[89]));
FA FA90 (.a(pp[8][15]),.b(pp[7][16]),.cin(pp[6][17]),.sum(fsu[90]),.carry(fca[90]));
FA FA91 (.a(pp[5][18]),.b(pp[4][19]),.cin(pp[3][20]),.sum(fsu[91]),.carry(fca[91]));
FA FA92 (.a(pp[2][21]),.b(pp[1][22]),.cin(pp[0][23]),.sum(fsu[92]),.carry(fca[92]));
FA FA93 (.a(pp[24][0]),.b(pp[23][1]),.cin(pp[22][2]),.sum(fsu[93]),.carry(fca[93]));
FA FA94 (.a(pp[21][3]),.b(pp[20][4]),.cin(pp[19][5]),.sum(fsu[94]),.carry(fca[94]));
FA FA95 (.a(pp[18][6]),.b(pp[17][7]),.cin(pp[16][8]),.sum(fsu[95]),.carry(fca[95]));
FA FA96 (.a(pp[15][9]),.b(pp[14][10]),.cin(pp[13][11]),.sum(fsu[96]),.carry(fca[96]));
FA FA97 (.a(pp[12][12]),.b(pp[11][13]),.cin(pp[10][14]),.sum(fsu[97]),.carry(fca[97]));
FA FA98 (.a(pp[9][15]),.b(pp[8][16]),.cin(pp[7][17]),.sum(fsu[98]),.carry(fca[98]));
FA FA99 (.a(pp[6][18]),.b(pp[5][19]),.cin(pp[4][20]),.sum(fsu[99]),.carry(fca[99]));
FA FA100 (.a(pp[3][21]),.b(pp[2][22]),.cin(pp[1][23]),.sum(fsu[100]),.carry(fca[100]));
FA FA101 (.a(pp[25][0]),.b(pp[24][1]),.cin(pp[23][2]),.sum(fsu[101]),.carry(fca[101]));
FA FA102 (.a(pp[22][3]),.b(pp[21][4]),.cin(pp[20][5]),.sum(fsu[102]),.carry(fca[102]));
FA FA103 (.a(pp[19][6]),.b(pp[18][7]),.cin(pp[17][8]),.sum(fsu[103]),.carry(fca[103]));
FA FA104 (.a(pp[16][9]),.b(pp[15][10]),.cin(pp[14][11]),.sum(fsu[104]),.carry(fca[104]));
FA FA105 (.a(pp[13][12]),.b(pp[12][13]),.cin(pp[11][14]),.sum(fsu[105]),.carry(fca[105]));
FA FA106 (.a(pp[10][15]),.b(pp[9][16]),.cin(pp[8][17]),.sum(fsu[106]),.carry(fca[106]));
FA FA107 (.a(pp[7][18]),.b(pp[6][19]),.cin(pp[5][20]),.sum(fsu[107]),.carry(fca[107]));
FA FA108 (.a(pp[4][21]),.b(pp[3][22]),.cin(pp[2][23]),.sum(fsu[108]),.carry(fca[108]));
HA HA9 (.a(pp[1][24]),.b(pp[0][25]),.sum_h(hsu[9]),.carry_h(hca[9]));
FA FA109 (.a(pp[26][0]),.b(pp[25][1]),.cin(pp[24][2]),.sum(fsu[109]),.carry(fca[109]));
FA FA110 (.a(pp[23][3]),.b(pp[22][4]),.cin(pp[21][5]),.sum(fsu[110]),.carry(fca[110]));
FA FA111 (.a(pp[20][6]),.b(pp[19][7]),.cin(pp[18][8]),.sum(fsu[111]),.carry(fca[111]));
FA FA112 (.a(pp[17][9]),.b(pp[16][10]),.cin(pp[15][11]),.sum(fsu[112]),.carry(fca[112]));
FA FA113 (.a(pp[14][12]),.b(pp[13][13]),.cin(pp[12][14]),.sum(fsu[113]),.carry(fca[113]));
FA FA114 (.a(pp[11][15]),.b(pp[10][16]),.cin(pp[9][17]),.sum(fsu[114]),.carry(fca[114]));
FA FA115 (.a(pp[8][18]),.b(pp[7][19]),.cin(pp[6][20]),.sum(fsu[115]),.carry(fca[115]));
FA FA116 (.a(pp[5][21]),.b(pp[4][22]),.cin(pp[3][23]),.sum(fsu[116]),.carry(fca[116]));
FA FA117 (.a(pp[2][24]),.b(pp[1][25]),.cin(pp[0][26]),.sum(fsu[117]),.carry(fca[117]));
FA FA118 (.a(pp[27][0]),.b(pp[26][1]),.cin(pp[25][2]),.sum(fsu[118]),.carry(fca[118]));
FA FA119 (.a(pp[24][3]),.b(pp[23][4]),.cin(pp[22][5]),.sum(fsu[119]),.carry(fca[119]));
FA FA120 (.a(pp[21][6]),.b(pp[20][7]),.cin(pp[19][8]),.sum(fsu[120]),.carry(fca[120]));
FA FA121 (.a(pp[18][9]),.b(pp[17][10]),.cin(pp[16][11]),.sum(fsu[121]),.carry(fca[121]));
FA FA122 (.a(pp[15][12]),.b(pp[14][13]),.cin(pp[13][14]),.sum(fsu[122]),.carry(fca[122]));
FA FA123 (.a(pp[12][15]),.b(pp[11][16]),.cin(pp[10][17]),.sum(fsu[123]),.carry(fca[123]));
FA FA124 (.a(pp[9][18]),.b(pp[8][19]),.cin(pp[7][20]),.sum(fsu[124]),.carry(fca[124]));
FA FA125 (.a(pp[6][21]),.b(pp[5][22]),.cin(pp[4][23]),.sum(fsu[125]),.carry(fca[125]));
FA FA126 (.a(pp[3][24]),.b(pp[2][25]),.cin(pp[1][26]),.sum(fsu[126]),.carry(fca[126]));
FA FA127 (.a(pp[28][0]),.b(pp[27][1]),.cin(pp[26][2]),.sum(fsu[127]),.carry(fca[127]));
FA FA128 (.a(pp[25][3]),.b(pp[24][4]),.cin(pp[23][5]),.sum(fsu[128]),.carry(fca[128]));
FA FA129 (.a(pp[22][6]),.b(pp[21][7]),.cin(pp[20][8]),.sum(fsu[129]),.carry(fca[129]));
FA FA130 (.a(pp[19][9]),.b(pp[18][10]),.cin(pp[17][11]),.sum(fsu[130]),.carry(fca[130]));
FA FA131 (.a(pp[16][12]),.b(pp[15][13]),.cin(pp[14][14]),.sum(fsu[131]),.carry(fca[131]));
FA FA132 (.a(pp[13][15]),.b(pp[12][16]),.cin(pp[11][17]),.sum(fsu[132]),.carry(fca[132]));
FA FA133 (.a(pp[10][18]),.b(pp[9][19]),.cin(pp[8][20]),.sum(fsu[133]),.carry(fca[133]));
FA FA134 (.a(pp[7][21]),.b(pp[6][22]),.cin(pp[5][23]),.sum(fsu[134]),.carry(fca[134]));
FA FA135 (.a(pp[4][24]),.b(pp[3][25]),.cin(pp[2][26]),.sum(fsu[135]),.carry(fca[135]));
HA HA10 (.a(pp[1][27]),.b(pp[0][28]),.sum_h(hsu[10]),.carry_h(hca[10]));
FA FA136 (.a(pp[29][0]),.b(pp[28][1]),.cin(pp[27][2]),.sum(fsu[136]),.carry(fca[136]));
FA FA137 (.a(pp[26][3]),.b(pp[25][4]),.cin(pp[24][5]),.sum(fsu[137]),.carry(fca[137]));
FA FA138 (.a(pp[23][6]),.b(pp[22][7]),.cin(pp[21][8]),.sum(fsu[138]),.carry(fca[138]));
FA FA139 (.a(pp[20][9]),.b(pp[19][10]),.cin(pp[18][11]),.sum(fsu[139]),.carry(fca[139]));
FA FA140 (.a(pp[17][12]),.b(pp[16][13]),.cin(pp[15][14]),.sum(fsu[140]),.carry(fca[140]));
FA FA141 (.a(pp[14][15]),.b(pp[13][16]),.cin(pp[12][17]),.sum(fsu[141]),.carry(fca[141]));
FA FA142 (.a(pp[11][18]),.b(pp[10][19]),.cin(pp[9][20]),.sum(fsu[142]),.carry(fca[142]));
FA FA143 (.a(pp[8][21]),.b(pp[7][22]),.cin(pp[6][23]),.sum(fsu[143]),.carry(fca[143]));
FA FA144 (.a(pp[5][24]),.b(pp[4][25]),.cin(pp[3][26]),.sum(fsu[144]),.carry(fca[144]));
FA FA145 (.a(pp[2][27]),.b(pp[1][28]),.cin(pp[0][29]),.sum(fsu[145]),.carry(fca[145]));
FA FA146 (.a(pp[30][0]),.b(pp[29][1]),.cin(pp[28][2]),.sum(fsu[146]),.carry(fca[146]));
FA FA147 (.a(pp[27][3]),.b(pp[26][4]),.cin(pp[25][5]),.sum(fsu[147]),.carry(fca[147]));
FA FA148 (.a(pp[24][6]),.b(pp[23][7]),.cin(pp[22][8]),.sum(fsu[148]),.carry(fca[148]));
FA FA149 (.a(pp[21][9]),.b(pp[20][10]),.cin(pp[19][11]),.sum(fsu[149]),.carry(fca[149]));
FA FA150 (.a(pp[18][12]),.b(pp[17][13]),.cin(pp[16][14]),.sum(fsu[150]),.carry(fca[150]));
FA FA151 (.a(pp[15][15]),.b(pp[14][16]),.cin(pp[13][17]),.sum(fsu[151]),.carry(fca[151]));
FA FA152 (.a(pp[12][18]),.b(pp[11][19]),.cin(pp[10][20]),.sum(fsu[152]),.carry(fca[152]));
FA FA153 (.a(pp[9][21]),.b(pp[8][22]),.cin(pp[7][23]),.sum(fsu[153]),.carry(fca[153]));
FA FA154 (.a(pp[6][24]),.b(pp[5][25]),.cin(pp[4][26]),.sum(fsu[154]),.carry(fca[154]));
FA FA155 (.a(pp[3][27]),.b(pp[2][28]),.cin(pp[1][29]),.sum(fsu[155]),.carry(fca[155]));
FA FA156 (.a(pp[31][0]),.b(pp[30][1]),.cin(pp[29][2]),.sum(fsu[156]),.carry(fca[156]));
FA FA157 (.a(pp[28][3]),.b(pp[27][4]),.cin(pp[26][5]),.sum(fsu[157]),.carry(fca[157]));
FA FA158 (.a(pp[25][6]),.b(pp[24][7]),.cin(pp[23][8]),.sum(fsu[158]),.carry(fca[158]));
FA FA159 (.a(pp[22][9]),.b(pp[21][10]),.cin(pp[20][11]),.sum(fsu[159]),.carry(fca[159]));
FA FA160 (.a(pp[19][12]),.b(pp[18][13]),.cin(pp[17][14]),.sum(fsu[160]),.carry(fca[160]));
FA FA161 (.a(pp[16][15]),.b(pp[15][16]),.cin(pp[14][17]),.sum(fsu[161]),.carry(fca[161]));
FA FA162 (.a(pp[13][18]),.b(pp[12][19]),.cin(pp[11][20]),.sum(fsu[162]),.carry(fca[162]));
FA FA163 (.a(pp[10][21]),.b(pp[9][22]),.cin(pp[8][23]),.sum(fsu[163]),.carry(fca[163]));
FA FA164 (.a(pp[7][24]),.b(pp[6][25]),.cin(pp[5][26]),.sum(fsu[164]),.carry(fca[164]));
FA FA165 (.a(pp[4][27]),.b(pp[3][28]),.cin(pp[2][29]),.sum(fsu[165]),.carry(fca[165]));
HA HA11 (.a(pp[31][1]),.b(pp[30][2]),.sum_h(hsu[11]),.carry_h(hca[11]));
FA FA166 (.a(pp[29][3]),.b(pp[28][4]),.cin(pp[27][5]),.sum(fsu[166]),.carry(fca[166]));
FA FA167 (.a(pp[26][6]),.b(pp[25][7]),.cin(pp[24][8]),.sum(fsu[167]),.carry(fca[167]));
FA FA168 (.a(pp[23][9]),.b(pp[22][10]),.cin(pp[21][11]),.sum(fsu[168]),.carry(fca[168]));
FA FA169 (.a(pp[20][12]),.b(pp[19][13]),.cin(pp[18][14]),.sum(fsu[169]),.carry(fca[169]));
FA FA170 (.a(pp[17][15]),.b(pp[16][16]),.cin(pp[15][17]),.sum(fsu[170]),.carry(fca[170]));
FA FA171 (.a(pp[14][18]),.b(pp[13][19]),.cin(pp[12][20]),.sum(fsu[171]),.carry(fca[171]));
FA FA172 (.a(pp[11][21]),.b(pp[10][22]),.cin(pp[9][23]),.sum(fsu[172]),.carry(fca[172]));
FA FA173 (.a(pp[8][24]),.b(pp[7][25]),.cin(pp[6][26]),.sum(fsu[173]),.carry(fca[173]));
FA FA174 (.a(pp[5][27]),.b(pp[4][28]),.cin(pp[3][29]),.sum(fsu[174]),.carry(fca[174]));
FA FA175 (.a(pp[30][3]),.b(pp[29][4]),.cin(pp[28][5]),.sum(fsu[175]),.carry(fca[175]));
FA FA176 (.a(pp[27][6]),.b(pp[26][7]),.cin(pp[25][8]),.sum(fsu[176]),.carry(fca[176]));
FA FA177 (.a(pp[24][9]),.b(pp[23][10]),.cin(pp[22][11]),.sum(fsu[177]),.carry(fca[177]));
FA FA178 (.a(pp[21][12]),.b(pp[20][13]),.cin(pp[19][14]),.sum(fsu[178]),.carry(fca[178]));
FA FA179 (.a(pp[18][15]),.b(pp[17][16]),.cin(pp[16][17]),.sum(fsu[179]),.carry(fca[179]));
FA FA180 (.a(pp[15][18]),.b(pp[14][19]),.cin(pp[13][20]),.sum(fsu[180]),.carry(fca[180]));
FA FA181 (.a(pp[12][21]),.b(pp[11][22]),.cin(pp[10][23]),.sum(fsu[181]),.carry(fca[181]));
FA FA182 (.a(pp[9][24]),.b(pp[8][25]),.cin(pp[7][26]),.sum(fsu[182]),.carry(fca[182]));
FA FA183 (.a(pp[6][27]),.b(pp[5][28]),.cin(pp[4][29]),.sum(fsu[183]),.carry(fca[183]));
FA FA184 (.a(pp[31][3]),.b(pp[30][4]),.cin(pp[29][5]),.sum(fsu[184]),.carry(fca[184]));
FA FA185 (.a(pp[28][6]),.b(pp[27][7]),.cin(pp[26][8]),.sum(fsu[185]),.carry(fca[185]));
FA FA186 (.a(pp[25][9]),.b(pp[24][10]),.cin(pp[23][11]),.sum(fsu[186]),.carry(fca[186]));
FA FA187 (.a(pp[22][12]),.b(pp[21][13]),.cin(pp[20][14]),.sum(fsu[187]),.carry(fca[187]));
FA FA188 (.a(pp[19][15]),.b(pp[18][16]),.cin(pp[17][17]),.sum(fsu[188]),.carry(fca[188]));
FA FA189 (.a(pp[16][18]),.b(pp[15][19]),.cin(pp[14][20]),.sum(fsu[189]),.carry(fca[189]));
FA FA190 (.a(pp[13][21]),.b(pp[12][22]),.cin(pp[11][23]),.sum(fsu[190]),.carry(fca[190]));
FA FA191 (.a(pp[10][24]),.b(pp[9][25]),.cin(pp[8][26]),.sum(fsu[191]),.carry(fca[191]));
FA FA192 (.a(pp[7][27]),.b(pp[6][28]),.cin(pp[5][29]),.sum(fsu[192]),.carry(fca[192]));
HA HA12 (.a(pp[31][4]),.b(pp[30][5]),.sum_h(hsu[12]),.carry_h(hca[12]));
FA FA193 (.a(pp[29][6]),.b(pp[28][7]),.cin(pp[27][8]),.sum(fsu[193]),.carry(fca[193]));
FA FA194 (.a(pp[26][9]),.b(pp[25][10]),.cin(pp[24][11]),.sum(fsu[194]),.carry(fca[194]));
FA FA195 (.a(pp[23][12]),.b(pp[22][13]),.cin(pp[21][14]),.sum(fsu[195]),.carry(fca[195]));
FA FA196 (.a(pp[20][15]),.b(pp[19][16]),.cin(pp[18][17]),.sum(fsu[196]),.carry(fca[196]));
FA FA197 (.a(pp[17][18]),.b(pp[16][19]),.cin(pp[15][20]),.sum(fsu[197]),.carry(fca[197]));
FA FA198 (.a(pp[14][21]),.b(pp[13][22]),.cin(pp[12][23]),.sum(fsu[198]),.carry(fca[198]));
FA FA199 (.a(pp[11][24]),.b(pp[10][25]),.cin(pp[9][26]),.sum(fsu[199]),.carry(fca[199]));
FA FA200 (.a(pp[8][27]),.b(pp[7][28]),.cin(pp[6][29]),.sum(fsu[200]),.carry(fca[200]));
FA FA201 (.a(pp[30][6]),.b(pp[29][7]),.cin(pp[28][8]),.sum(fsu[201]),.carry(fca[201]));
FA FA202 (.a(pp[27][9]),.b(pp[26][10]),.cin(pp[25][11]),.sum(fsu[202]),.carry(fca[202]));
FA FA203 (.a(pp[24][12]),.b(pp[23][13]),.cin(pp[22][14]),.sum(fsu[203]),.carry(fca[203]));
FA FA204 (.a(pp[21][15]),.b(pp[20][16]),.cin(pp[19][17]),.sum(fsu[204]),.carry(fca[204]));
FA FA205 (.a(pp[18][18]),.b(pp[17][19]),.cin(pp[16][20]),.sum(fsu[205]),.carry(fca[205]));
FA FA206 (.a(pp[15][21]),.b(pp[14][22]),.cin(pp[13][23]),.sum(fsu[206]),.carry(fca[206]));
FA FA207 (.a(pp[12][24]),.b(pp[11][25]),.cin(pp[10][26]),.sum(fsu[207]),.carry(fca[207]));
FA FA208 (.a(pp[9][27]),.b(pp[8][28]),.cin(pp[7][29]),.sum(fsu[208]),.carry(fca[208]));
FA FA209 (.a(pp[31][6]),.b(pp[30][7]),.cin(pp[29][8]),.sum(fsu[209]),.carry(fca[209]));
FA FA210 (.a(pp[28][9]),.b(pp[27][10]),.cin(pp[26][11]),.sum(fsu[210]),.carry(fca[210]));
FA FA211 (.a(pp[25][12]),.b(pp[24][13]),.cin(pp[23][14]),.sum(fsu[211]),.carry(fca[211]));
FA FA212 (.a(pp[22][15]),.b(pp[21][16]),.cin(pp[20][17]),.sum(fsu[212]),.carry(fca[212]));
FA FA213 (.a(pp[19][18]),.b(pp[18][19]),.cin(pp[17][20]),.sum(fsu[213]),.carry(fca[213]));
FA FA214 (.a(pp[16][21]),.b(pp[15][22]),.cin(pp[14][23]),.sum(fsu[214]),.carry(fca[214]));
FA FA215 (.a(pp[13][24]),.b(pp[12][25]),.cin(pp[11][26]),.sum(fsu[215]),.carry(fca[215]));
FA FA216 (.a(pp[10][27]),.b(pp[9][28]),.cin(pp[8][29]),.sum(fsu[216]),.carry(fca[216]));
HA HA13 (.a(pp[31][7]),.b(pp[30][8]),.sum_h(hsu[13]),.carry_h(hca[13]));
FA FA217 (.a(pp[29][9]),.b(pp[28][10]),.cin(pp[27][11]),.sum(fsu[217]),.carry(fca[217]));
FA FA218 (.a(pp[26][12]),.b(pp[25][13]),.cin(pp[24][14]),.sum(fsu[218]),.carry(fca[218]));
FA FA219 (.a(pp[23][15]),.b(pp[22][16]),.cin(pp[21][17]),.sum(fsu[219]),.carry(fca[219]));
FA FA220 (.a(pp[20][18]),.b(pp[19][19]),.cin(pp[18][20]),.sum(fsu[220]),.carry(fca[220]));
FA FA221 (.a(pp[17][21]),.b(pp[16][22]),.cin(pp[15][23]),.sum(fsu[221]),.carry(fca[221]));
FA FA222 (.a(pp[14][24]),.b(pp[13][25]),.cin(pp[12][26]),.sum(fsu[222]),.carry(fca[222]));
FA FA223 (.a(pp[11][27]),.b(pp[10][28]),.cin(pp[9][29]),.sum(fsu[223]),.carry(fca[223]));
FA FA224 (.a(pp[30][9]),.b(pp[29][10]),.cin(pp[28][11]),.sum(fsu[224]),.carry(fca[224]));
FA FA225 (.a(pp[27][12]),.b(pp[26][13]),.cin(pp[25][14]),.sum(fsu[225]),.carry(fca[225]));
FA FA226 (.a(pp[24][15]),.b(pp[23][16]),.cin(pp[22][17]),.sum(fsu[226]),.carry(fca[226]));
FA FA227 (.a(pp[21][18]),.b(pp[20][19]),.cin(pp[19][20]),.sum(fsu[227]),.carry(fca[227]));
FA FA228 (.a(pp[18][21]),.b(pp[17][22]),.cin(pp[16][23]),.sum(fsu[228]),.carry(fca[228]));
FA FA229 (.a(pp[15][24]),.b(pp[14][25]),.cin(pp[13][26]),.sum(fsu[229]),.carry(fca[229]));
FA FA230 (.a(pp[12][27]),.b(pp[11][28]),.cin(pp[10][29]),.sum(fsu[230]),.carry(fca[230]));
FA FA231 (.a(pp[31][9]),.b(pp[30][10]),.cin(pp[29][11]),.sum(fsu[231]),.carry(fca[231]));
FA FA232 (.a(pp[28][12]),.b(pp[27][13]),.cin(pp[26][14]),.sum(fsu[232]),.carry(fca[232]));
FA FA233 (.a(pp[25][15]),.b(pp[24][16]),.cin(pp[23][17]),.sum(fsu[233]),.carry(fca[233]));
FA FA234 (.a(pp[22][18]),.b(pp[21][19]),.cin(pp[20][20]),.sum(fsu[234]),.carry(fca[234]));
FA FA235 (.a(pp[19][21]),.b(pp[18][22]),.cin(pp[17][23]),.sum(fsu[235]),.carry(fca[235]));
FA FA236 (.a(pp[16][24]),.b(pp[15][25]),.cin(pp[14][26]),.sum(fsu[236]),.carry(fca[236]));
FA FA237 (.a(pp[13][27]),.b(pp[12][28]),.cin(pp[11][29]),.sum(fsu[237]),.carry(fca[237]));
HA HA14 (.a(pp[31][10]),.b(pp[30][11]),.sum_h(hsu[14]),.carry_h(hca[14]));
FA FA238 (.a(pp[29][12]),.b(pp[28][13]),.cin(pp[27][14]),.sum(fsu[238]),.carry(fca[238]));
FA FA239 (.a(pp[26][15]),.b(pp[25][16]),.cin(pp[24][17]),.sum(fsu[239]),.carry(fca[239]));
FA FA240 (.a(pp[23][18]),.b(pp[22][19]),.cin(pp[21][20]),.sum(fsu[240]),.carry(fca[240]));
FA FA241 (.a(pp[20][21]),.b(pp[19][22]),.cin(pp[18][23]),.sum(fsu[241]),.carry(fca[241]));
FA FA242 (.a(pp[17][24]),.b(pp[16][25]),.cin(pp[15][26]),.sum(fsu[242]),.carry(fca[242]));
FA FA243 (.a(pp[14][27]),.b(pp[13][28]),.cin(pp[12][29]),.sum(fsu[243]),.carry(fca[243]));
FA FA244 (.a(pp[30][12]),.b(pp[29][13]),.cin(pp[28][14]),.sum(fsu[244]),.carry(fca[244]));
FA FA245 (.a(pp[27][15]),.b(pp[26][16]),.cin(pp[25][17]),.sum(fsu[245]),.carry(fca[245]));
FA FA246 (.a(pp[24][18]),.b(pp[23][19]),.cin(pp[22][20]),.sum(fsu[246]),.carry(fca[246]));
FA FA247 (.a(pp[21][21]),.b(pp[20][22]),.cin(pp[19][23]),.sum(fsu[247]),.carry(fca[247]));
FA FA248 (.a(pp[18][24]),.b(pp[17][25]),.cin(pp[16][26]),.sum(fsu[248]),.carry(fca[248]));
FA FA249 (.a(pp[15][27]),.b(pp[14][28]),.cin(pp[13][29]),.sum(fsu[249]),.carry(fca[249]));
FA FA250 (.a(pp[31][12]),.b(pp[30][13]),.cin(pp[29][14]),.sum(fsu[250]),.carry(fca[250]));
FA FA251 (.a(pp[28][15]),.b(pp[27][16]),.cin(pp[26][17]),.sum(fsu[251]),.carry(fca[251]));
FA FA252 (.a(pp[25][18]),.b(pp[24][19]),.cin(pp[23][20]),.sum(fsu[252]),.carry(fca[252]));
FA FA253 (.a(pp[22][21]),.b(pp[21][22]),.cin(pp[20][23]),.sum(fsu[253]),.carry(fca[253]));
FA FA254 (.a(pp[19][24]),.b(pp[18][25]),.cin(pp[17][26]),.sum(fsu[254]),.carry(fca[254]));
FA FA255 (.a(pp[16][27]),.b(pp[15][28]),.cin(pp[14][29]),.sum(fsu[255]),.carry(fca[255]));
HA HA15 (.a(pp[31][13]),.b(pp[30][14]),.sum_h(hsu[15]),.carry_h(hca[15]));
FA FA256 (.a(pp[29][15]),.b(pp[28][16]),.cin(pp[27][17]),.sum(fsu[256]),.carry(fca[256]));
FA FA257 (.a(pp[26][18]),.b(pp[25][19]),.cin(pp[24][20]),.sum(fsu[257]),.carry(fca[257]));
FA FA258 (.a(pp[23][21]),.b(pp[22][22]),.cin(pp[21][23]),.sum(fsu[258]),.carry(fca[258]));
FA FA259 (.a(pp[20][24]),.b(pp[19][25]),.cin(pp[18][26]),.sum(fsu[259]),.carry(fca[259]));
FA FA260 (.a(pp[17][27]),.b(pp[16][28]),.cin(pp[15][29]),.sum(fsu[260]),.carry(fca[260]));
FA FA261 (.a(pp[30][15]),.b(pp[29][16]),.cin(pp[28][17]),.sum(fsu[261]),.carry(fca[261]));
FA FA262 (.a(pp[27][18]),.b(pp[26][19]),.cin(pp[25][20]),.sum(fsu[262]),.carry(fca[262]));
FA FA263 (.a(pp[24][21]),.b(pp[23][22]),.cin(pp[22][23]),.sum(fsu[263]),.carry(fca[263]));
FA FA264 (.a(pp[21][24]),.b(pp[20][25]),.cin(pp[19][26]),.sum(fsu[264]),.carry(fca[264]));
FA FA265 (.a(pp[18][27]),.b(pp[17][28]),.cin(pp[16][29]),.sum(fsu[265]),.carry(fca[265]));
FA FA266 (.a(pp[31][15]),.b(pp[30][16]),.cin(pp[29][17]),.sum(fsu[266]),.carry(fca[266]));
FA FA267 (.a(pp[28][18]),.b(pp[27][19]),.cin(pp[26][20]),.sum(fsu[267]),.carry(fca[267]));
FA FA268 (.a(pp[25][21]),.b(pp[24][22]),.cin(pp[23][23]),.sum(fsu[268]),.carry(fca[268]));
FA FA269 (.a(pp[22][24]),.b(pp[21][25]),.cin(pp[20][26]),.sum(fsu[269]),.carry(fca[269]));
FA FA270 (.a(pp[19][27]),.b(pp[18][28]),.cin(pp[17][29]),.sum(fsu[270]),.carry(fca[270]));
HA HA16 (.a(pp[31][16]),.b(pp[30][17]),.sum_h(hsu[16]),.carry_h(hca[16]));
FA FA271 (.a(pp[29][18]),.b(pp[28][19]),.cin(pp[27][20]),.sum(fsu[271]),.carry(fca[271]));
FA FA272 (.a(pp[26][21]),.b(pp[25][22]),.cin(pp[24][23]),.sum(fsu[272]),.carry(fca[272]));
FA FA273 (.a(pp[23][24]),.b(pp[22][25]),.cin(pp[21][26]),.sum(fsu[273]),.carry(fca[273]));
FA FA274 (.a(pp[20][27]),.b(pp[19][28]),.cin(pp[18][29]),.sum(fsu[274]),.carry(fca[274]));
FA FA275 (.a(pp[30][18]),.b(pp[29][19]),.cin(pp[28][20]),.sum(fsu[275]),.carry(fca[275]));
FA FA276 (.a(pp[27][21]),.b(pp[26][22]),.cin(pp[25][23]),.sum(fsu[276]),.carry(fca[276]));
FA FA277 (.a(pp[24][24]),.b(pp[23][25]),.cin(pp[22][26]),.sum(fsu[277]),.carry(fca[277]));
FA FA278 (.a(pp[21][27]),.b(pp[20][28]),.cin(pp[19][29]),.sum(fsu[278]),.carry(fca[278]));
FA FA279 (.a(pp[31][18]),.b(pp[30][19]),.cin(pp[29][20]),.sum(fsu[279]),.carry(fca[279]));
FA FA280 (.a(pp[28][21]),.b(pp[27][22]),.cin(pp[26][23]),.sum(fsu[280]),.carry(fca[280]));
FA FA281 (.a(pp[25][24]),.b(pp[24][25]),.cin(pp[23][26]),.sum(fsu[281]),.carry(fca[281]));
FA FA282 (.a(pp[22][27]),.b(pp[21][28]),.cin(pp[20][29]),.sum(fsu[282]),.carry(fca[282]));
HA HA17 (.a(pp[31][19]),.b(pp[30][20]),.sum_h(hsu[17]),.carry_h(hca[17]));
FA FA283 (.a(pp[29][21]),.b(pp[28][22]),.cin(pp[27][23]),.sum(fsu[283]),.carry(fca[283]));
FA FA284 (.a(pp[26][24]),.b(pp[25][25]),.cin(pp[24][26]),.sum(fsu[284]),.carry(fca[284]));
FA FA285 (.a(pp[23][27]),.b(pp[22][28]),.cin(pp[21][29]),.sum(fsu[285]),.carry(fca[285]));
FA FA286 (.a(pp[30][21]),.b(pp[29][22]),.cin(pp[28][23]),.sum(fsu[286]),.carry(fca[286]));
FA FA287 (.a(pp[27][24]),.b(pp[26][25]),.cin(pp[25][26]),.sum(fsu[287]),.carry(fca[287]));
FA FA288 (.a(pp[24][27]),.b(pp[23][28]),.cin(pp[22][29]),.sum(fsu[288]),.carry(fca[288]));
FA FA289 (.a(pp[31][21]),.b(pp[30][22]),.cin(pp[29][23]),.sum(fsu[289]),.carry(fca[289]));
FA FA290 (.a(pp[28][24]),.b(pp[27][25]),.cin(pp[26][26]),.sum(fsu[290]),.carry(fca[290]));
FA FA291 (.a(pp[25][27]),.b(pp[24][28]),.cin(pp[23][29]),.sum(fsu[291]),.carry(fca[291]));
HA HA18 (.a(pp[31][22]),.b(pp[30][23]),.sum_h(hsu[18]),.carry_h(hca[18]));
FA FA292 (.a(pp[29][24]),.b(pp[28][25]),.cin(pp[27][26]),.sum(fsu[292]),.carry(fca[292]));
FA FA293 (.a(pp[26][27]),.b(pp[25][28]),.cin(pp[24][29]),.sum(fsu[293]),.carry(fca[293]));
FA FA294 (.a(pp[30][24]),.b(pp[29][25]),.cin(pp[28][26]),.sum(fsu[294]),.carry(fca[294]));
FA FA295 (.a(pp[27][27]),.b(pp[26][28]),.cin(pp[25][29]),.sum(fsu[295]),.carry(fca[295]));
FA FA296 (.a(pp[31][24]),.b(pp[30][25]),.cin(pp[29][26]),.sum(fsu[296]),.carry(fca[296]));
FA FA297 (.a(pp[28][27]),.b(pp[27][28]),.cin(pp[26][29]),.sum(fsu[297]),.carry(fca[297]));
HA HA19 (.a(pp[31][25]),.b(pp[30][26]),.sum_h(hsu[19]),.carry_h(hca[19]));
FA FA298 (.a(pp[29][27]),.b(pp[28][28]),.cin(pp[27][29]),.sum(fsu[298]),.carry(fca[298]));
FA FA299 (.a(pp[30][27]),.b(pp[29][28]),.cin(pp[28][29]),.sum(fsu[299]),.carry(fca[299]));
FA FA300 (.a(pp[31][27]),.b(pp[30][28]),.cin(pp[29][29]),.sum(fsu[300]),.carry(fca[300]));
HA HA20 (.a(pp[31][28]),.b(pp[30][29]),.sum_h(hsu[20]),.carry_h(hca[20]));
//2nd stage
HA HA21 (.a(fsu[1]),.b(hca[1]),.sum_h(z[2]),.carry_h(hca[21]));
FA FA301 (.a(fsu[2]),.b(fca[1]),.cin(pp[0][3]),.sum(fsu[301]),.carry(fca[301]));
FA FA302 (.a(fsu[3]),.b(fca[2]),.cin(hsu[2]),.sum(fsu[302]),.carry(fca[302]));
FA FA303 (.a(fsu[4]),.b(fca[3]),.cin(fsu[5]),.sum(fsu[303]),.carry(fca[303]));
FA FA304 (.a(fsu[6]),.b(fca[4]),.cin(fsu[7]),.sum(fsu[304]),.carry(fca[304]));
HA HA22 (.a(fca[5]),.b(pp[0][6]),.sum_h(hsu[22]),.carry_h(hca[22]));
FA FA305 (.a(fsu[8]),.b(fca[6]),.cin(fsu[9]),.sum(fsu[305]),.carry(fca[305]));
HA HA23 (.a(fca[7]),.b(hsu[3]),.sum_h(hsu[23]),.carry_h(hca[23]));
FA FA306 (.a(fsu[10]),.b(fca[8]),.cin(fsu[11]),.sum(fsu[306]),.carry(fca[306]));
FA FA307 (.a(fca[9]),.b(fsu[12]),.cin(hca[3]),.sum(fsu[307]),.carry(fca[307]));
FA FA308 (.a(fsu[13]),.b(fca[10]),.cin(fsu[14]),.sum(fsu[308]),.carry(fca[308]));
FA FA309 (.a(fca[11]),.b(fsu[15]),.cin(fca[12]),.sum(fsu[309]),.carry(fca[309]));
FA FA310 (.a(fsu[16]),.b(fca[13]),.cin(fsu[17]),.sum(fsu[310]),.carry(fca[310]));
FA FA311 (.a(fca[14]),.b(fsu[18]),.cin(fca[15]),.sum(fsu[311]),.carry(fca[311]));
FA FA312 (.a(fsu[19]),.b(fca[16]),.cin(fsu[20]),.sum(fsu[312]),.carry(fca[312]));
FA FA313 (.a(fca[17]),.b(fsu[21]),.cin(fca[18]),.sum(fsu[313]),.carry(fca[313]));
HA HA24 (.a(fsu[22]),.b(hca[4]),.sum_h(hsu[24]),.carry_h(hca[24]));
FA FA314 (.a(fsu[23]),.b(fca[19]),.cin(fsu[24]),.sum(fsu[314]),.carry(fca[314]));
FA FA315 (.a(fca[20]),.b(fsu[25]),.cin(fca[21]),.sum(fsu[315]),.carry(fca[315]));
FA FA316 (.a(fsu[26]),.b(fca[22]),.cin(pp[0][12]),.sum(fsu[316]),.carry(fca[316]));
FA FA317 (.a(fsu[27]),.b(fca[23]),.cin(fsu[28]),.sum(fsu[317]),.carry(fca[317]));
FA FA318 (.a(fca[24]),.b(fsu[29]),.cin(fca[25]),.sum(fsu[318]),.carry(fca[318]));
FA FA319 (.a(fsu[30]),.b(fca[26]),.cin(hsu[5]),.sum(fsu[319]),.carry(fca[319]));
FA FA320 (.a(fsu[31]),.b(fca[27]),.cin(fsu[32]),.sum(fsu[320]),.carry(fca[320]));
FA FA321 (.a(fca[28]),.b(fsu[33]),.cin(fca[29]),.sum(fsu[321]),.carry(fca[321]));
FA FA322 (.a(fsu[34]),.b(fca[30]),.cin(fsu[35]),.sum(fsu[322]),.carry(fca[322]));
FA FA323 (.a(fsu[36]),.b(fca[31]),.cin(fsu[37]),.sum(fsu[323]),.carry(fca[323]));
FA FA324 (.a(fca[32]),.b(fsu[38]),.cin(fca[33]),.sum(fsu[324]),.carry(fca[324]));
FA FA325 (.a(fsu[39]),.b(fca[34]),.cin(fsu[40]),.sum(fsu[325]),.carry(fca[325]));
HA HA25 (.a(fca[35]),.b(pp[0][15]),.sum_h(hsu[25]),.carry_h(hca[25]));
FA FA326 (.a(fsu[41]),.b(fca[36]),.cin(fsu[42]),.sum(fsu[326]),.carry(fca[326]));
FA FA327 (.a(fca[37]),.b(fsu[43]),.cin(fca[38]),.sum(fsu[327]),.carry(fca[327]));
FA FA328 (.a(fsu[44]),.b(fca[39]),.cin(fsu[45]),.sum(fsu[328]),.carry(fca[328]));
HA HA26 (.a(fca[40]),.b(hsu[6]),.sum_h(hsu[26]),.carry_h(hca[26]));
FA FA329 (.a(fsu[46]),.b(fca[41]),.cin(fsu[47]),.sum(fsu[329]),.carry(fca[329]));
FA FA330 (.a(fca[42]),.b(fsu[48]),.cin(fca[43]),.sum(fsu[330]),.carry(fca[330]));
FA FA331 (.a(fsu[49]),.b(fca[44]),.cin(fsu[50]),.sum(fsu[331]),.carry(fca[331]));
FA FA332 (.a(fca[45]),.b(fsu[51]),.cin(hca[6]),.sum(fsu[332]),.carry(fca[332]));
FA FA333 (.a(fsu[52]),.b(fca[46]),.cin(fsu[53]),.sum(fsu[333]),.carry(fca[333]));
FA FA334 (.a(fca[47]),.b(fsu[54]),.cin(fca[48]),.sum(fsu[334]),.carry(fca[334]));
FA FA335 (.a(fsu[55]),.b(fca[49]),.cin(fsu[56]),.sum(fsu[335]),.carry(fca[335]));
FA FA336 (.a(fca[50]),.b(fsu[57]),.cin(fca[51]),.sum(fsu[336]),.carry(fca[336]));
FA FA337 (.a(fsu[58]),.b(fca[52]),.cin(fsu[59]),.sum(fsu[337]),.carry(fca[337]));
FA FA338 (.a(fca[53]),.b(fsu[60]),.cin(fca[54]),.sum(fsu[338]),.carry(fca[338]));
FA FA339 (.a(fsu[61]),.b(fca[55]),.cin(fsu[62]),.sum(fsu[339]),.carry(fca[339]));
FA FA340 (.a(fca[56]),.b(fsu[63]),.cin(fca[57]),.sum(fsu[340]),.carry(fca[340]));
FA FA341 (.a(fsu[64]),.b(fca[58]),.cin(fsu[65]),.sum(fsu[341]),.carry(fca[341]));
FA FA342 (.a(fca[59]),.b(fsu[66]),.cin(fca[60]),.sum(fsu[342]),.carry(fca[342]));
FA FA343 (.a(fsu[67]),.b(fca[61]),.cin(fsu[68]),.sum(fsu[343]),.carry(fca[343]));
FA FA344 (.a(fca[62]),.b(fsu[69]),.cin(fca[63]),.sum(fsu[344]),.carry(fca[344]));
HA HA27 (.a(fsu[70]),.b(hca[7]),.sum_h(hsu[27]),.carry_h(hca[27]));
FA FA345 (.a(fsu[71]),.b(fca[64]),.cin(fsu[72]),.sum(fsu[345]),.carry(fca[345]));
FA FA346 (.a(fca[65]),.b(fsu[73]),.cin(fca[66]),.sum(fsu[346]),.carry(fca[346]));
FA FA347 (.a(fsu[74]),.b(fca[67]),.cin(fsu[75]),.sum(fsu[347]),.carry(fca[347]));
FA FA348 (.a(fca[68]),.b(fsu[76]),.cin(fca[69]),.sum(fsu[348]),.carry(fca[348]));
FA FA349 (.a(fsu[77]),.b(fca[70]),.cin(pp[0][21]),.sum(fsu[349]),.carry(fca[349]));
FA FA350 (.a(fsu[78]),.b(fca[71]),.cin(fsu[79]),.sum(fsu[350]),.carry(fca[350]));
FA FA351 (.a(fca[72]),.b(fsu[80]),.cin(fca[73]),.sum(fsu[351]),.carry(fca[351]));
FA FA352 (.a(fsu[81]),.b(fca[74]),.cin(fsu[82]),.sum(fsu[352]),.carry(fca[352]));
FA FA353 (.a(fca[75]),.b(fsu[83]),.cin(fca[76]),.sum(fsu[353]),.carry(fca[353]));
FA FA354 (.a(fsu[84]),.b(fca[77]),.cin(hsu[8]),.sum(fsu[354]),.carry(fca[354]));
FA FA355 (.a(fsu[85]),.b(fca[78]),.cin(fsu[86]),.sum(fsu[355]),.carry(fca[355]));
FA FA356 (.a(fca[79]),.b(fsu[87]),.cin(fca[80]),.sum(fsu[356]),.carry(fca[356]));
FA FA357 (.a(fsu[88]),.b(fca[81]),.cin(fsu[89]),.sum(fsu[357]),.carry(fca[357]));
FA FA358 (.a(fca[82]),.b(fsu[90]),.cin(fca[83]),.sum(fsu[358]),.carry(fca[358]));
FA FA359 (.a(fsu[91]),.b(fca[84]),.cin(fsu[92]),.sum(fsu[359]),.carry(fca[359]));
FA FA360 (.a(fsu[93]),.b(fca[85]),.cin(fsu[94]),.sum(fsu[360]),.carry(fca[360]));
FA FA361 (.a(fca[86]),.b(fsu[95]),.cin(fca[87]),.sum(fsu[361]),.carry(fca[361]));
FA FA362 (.a(fsu[96]),.b(fca[88]),.cin(fsu[97]),.sum(fsu[362]),.carry(fca[362]));
FA FA363 (.a(fca[89]),.b(fsu[98]),.cin(fca[90]),.sum(fsu[363]),.carry(fca[363]));
FA FA364 (.a(fsu[99]),.b(fca[91]),.cin(fsu[100]),.sum(fsu[364]),.carry(fca[364]));
HA HA28 (.a(fca[92]),.b(pp[0][24]),.sum_h(hsu[28]),.carry_h(hca[28]));
FA FA365 (.a(fsu[101]),.b(fca[93]),.cin(fsu[102]),.sum(fsu[365]),.carry(fca[365]));
FA FA366 (.a(fca[94]),.b(fsu[103]),.cin(fca[95]),.sum(fsu[366]),.carry(fca[366]));
FA FA367 (.a(fsu[104]),.b(fca[96]),.cin(fsu[105]),.sum(fsu[367]),.carry(fca[367]));
FA FA368 (.a(fca[97]),.b(fsu[106]),.cin(fca[98]),.sum(fsu[368]),.carry(fca[368]));
FA FA369 (.a(fsu[107]),.b(fca[99]),.cin(fsu[108]),.sum(fsu[369]),.carry(fca[369]));
HA HA29 (.a(fca[100]),.b(hsu[9]),.sum_h(hsu[29]),.carry_h(hca[29]));
FA FA370 (.a(fsu[109]),.b(fca[101]),.cin(fsu[110]),.sum(fsu[370]),.carry(fca[370]));
FA FA371 (.a(fca[102]),.b(fsu[111]),.cin(fca[103]),.sum(fsu[371]),.carry(fca[371]));
FA FA372 (.a(fsu[112]),.b(fca[104]),.cin(fsu[113]),.sum(fsu[372]),.carry(fca[372]));
FA FA373 (.a(fca[105]),.b(fsu[114]),.cin(fca[106]),.sum(fsu[373]),.carry(fca[373]));
FA FA374 (.a(fsu[115]),.b(fca[107]),.cin(fsu[116]),.sum(fsu[374]),.carry(fca[374]));
FA FA375 (.a(fca[108]),.b(fsu[117]),.cin(hca[9]),.sum(fsu[375]),.carry(fca[375]));
FA FA376 (.a(fsu[118]),.b(fca[109]),.cin(fsu[119]),.sum(fsu[376]),.carry(fca[376]));
FA FA377 (.a(fca[110]),.b(fsu[120]),.cin(fca[111]),.sum(fsu[377]),.carry(fca[377]));
FA FA378 (.a(fsu[121]),.b(fca[112]),.cin(fsu[122]),.sum(fsu[378]),.carry(fca[378]));
FA FA379 (.a(fca[113]),.b(fsu[123]),.cin(fca[114]),.sum(fsu[379]),.carry(fca[379]));
FA FA380 (.a(fsu[124]),.b(fca[115]),.cin(fsu[125]),.sum(fsu[380]),.carry(fca[380]));
FA FA381 (.a(fca[116]),.b(fsu[126]),.cin(fca[117]),.sum(fsu[381]),.carry(fca[381]));
FA FA382 (.a(fsu[127]),.b(fca[118]),.cin(fsu[128]),.sum(fsu[382]),.carry(fca[382]));
FA FA383 (.a(fca[119]),.b(fsu[129]),.cin(fca[120]),.sum(fsu[383]),.carry(fca[383]));
FA FA384 (.a(fsu[130]),.b(fca[121]),.cin(fsu[131]),.sum(fsu[384]),.carry(fca[384]));
FA FA385 (.a(fca[122]),.b(fsu[132]),.cin(fca[123]),.sum(fsu[385]),.carry(fca[385]));
FA FA386 (.a(fsu[133]),.b(fca[124]),.cin(fsu[134]),.sum(fsu[386]),.carry(fca[386]));
FA FA387 (.a(fca[125]),.b(fsu[135]),.cin(fca[126]),.sum(fsu[387]),.carry(fca[387]));
FA FA388 (.a(fsu[136]),.b(fca[127]),.cin(fsu[137]),.sum(fsu[388]),.carry(fca[388]));
FA FA389 (.a(fca[128]),.b(fsu[138]),.cin(fca[129]),.sum(fsu[389]),.carry(fca[389]));
FA FA390 (.a(fsu[139]),.b(fca[130]),.cin(fsu[140]),.sum(fsu[390]),.carry(fca[390]));
FA FA391 (.a(fca[131]),.b(fsu[141]),.cin(fca[132]),.sum(fsu[391]),.carry(fca[391]));
FA FA392 (.a(fsu[142]),.b(fca[133]),.cin(fsu[143]),.sum(fsu[392]),.carry(fca[392]));
FA FA393 (.a(fca[134]),.b(fsu[144]),.cin(fca[135]),.sum(fsu[393]),.carry(fca[393]));
HA HA30 (.a(fsu[145]),.b(hca[10]),.sum_h(hsu[30]),.carry_h(hca[30]));
FA FA394 (.a(fsu[146]),.b(fca[136]),.cin(fsu[147]),.sum(fsu[394]),.carry(fca[394]));
FA FA395 (.a(fca[137]),.b(fsu[148]),.cin(fca[138]),.sum(fsu[395]),.carry(fca[395]));
FA FA396 (.a(fsu[149]),.b(fca[139]),.cin(fsu[150]),.sum(fsu[396]),.carry(fca[396]));
FA FA397 (.a(fca[140]),.b(fsu[151]),.cin(fca[141]),.sum(fsu[397]),.carry(fca[397]));
FA FA398 (.a(fsu[152]),.b(fca[142]),.cin(fsu[153]),.sum(fsu[398]),.carry(fca[398]));
FA FA399 (.a(fca[143]),.b(fsu[154]),.cin(fca[144]),.sum(fsu[399]),.carry(fca[399]));
FA FA400 (.a(fsu[155]),.b(fca[145]),.cin(pp[0][30]),.sum(fsu[400]),.carry(fca[400]));
FA FA401 (.a(fsu[156]),.b(fca[146]),.cin(fsu[157]),.sum(fsu[401]),.carry(fca[401]));
FA FA402 (.a(fca[147]),.b(fsu[158]),.cin(fca[148]),.sum(fsu[402]),.carry(fca[402]));
FA FA403 (.a(fsu[159]),.b(fca[149]),.cin(fsu[160]),.sum(fsu[403]),.carry(fca[403]));
FA FA404 (.a(fca[150]),.b(fsu[161]),.cin(fca[151]),.sum(fsu[404]),.carry(fca[404]));
FA FA405 (.a(fsu[162]),.b(fca[152]),.cin(fsu[163]),.sum(fsu[405]),.carry(fca[405]));
FA FA406 (.a(fca[153]),.b(fsu[164]),.cin(fca[154]),.sum(fsu[406]),.carry(fca[406]));
FA FA407 (.a(fsu[165]),.b(fca[155]),.cin(pp[1][30]),.sum(fsu[407]),.carry(fca[407]));
FA FA408 (.a(hsu[11]),.b(fca[156]),.cin(fsu[166]),.sum(fsu[408]),.carry(fca[408]));
FA FA409 (.a(fca[157]),.b(fsu[167]),.cin(fca[158]),.sum(fsu[409]),.carry(fca[409]));
FA FA410 (.a(fsu[168]),.b(fca[159]),.cin(fsu[169]),.sum(fsu[410]),.carry(fca[410]));
FA FA411 (.a(fca[160]),.b(fsu[170]),.cin(fca[161]),.sum(fsu[411]),.carry(fca[411]));
FA FA412 (.a(fsu[171]),.b(fca[162]),.cin(fsu[172]),.sum(fsu[412]),.carry(fca[412]));
FA FA413 (.a(fca[163]),.b(fsu[173]),.cin(fca[164]),.sum(fsu[413]),.carry(fca[413]));
FA FA414 (.a(fsu[174]),.b(fca[165]),.cin(pp[2][30]),.sum(fsu[414]),.carry(fca[414]));
FA FA415 (.a(pp[31][2]),.b(hca[11]),.cin(fsu[175]),.sum(fsu[415]),.carry(fca[415]));
FA FA416 (.a(fca[166]),.b(fsu[176]),.cin(fca[167]),.sum(fsu[416]),.carry(fca[416]));
FA FA417 (.a(fsu[177]),.b(fca[168]),.cin(fsu[178]),.sum(fsu[417]),.carry(fca[417]));
FA FA418 (.a(fca[169]),.b(fsu[179]),.cin(fca[170]),.sum(fsu[418]),.carry(fca[418]));
FA FA419 (.a(fsu[180]),.b(fca[171]),.cin(fsu[181]),.sum(fsu[419]),.carry(fca[419]));
FA FA420 (.a(fca[172]),.b(fsu[182]),.cin(fca[173]),.sum(fsu[420]),.carry(fca[420]));
FA FA421 (.a(fsu[183]),.b(fca[174]),.cin(pp[3][30]),.sum(fsu[421]),.carry(fca[421]));
FA FA422 (.a(fca[175]),.b(fsu[185]),.cin(fca[176]),.sum(fsu[422]),.carry(fca[422]));
FA FA423 (.a(fsu[186]),.b(fca[177]),.cin(fsu[187]),.sum(fsu[423]),.carry(fca[423]));
FA FA424 (.a(fca[178]),.b(fsu[188]),.cin(fca[179]),.sum(fsu[424]),.carry(fca[424]));
FA FA425 (.a(fsu[189]),.b(fca[180]),.cin(fsu[190]),.sum(fsu[425]),.carry(fca[425]));
FA FA426 (.a(fca[181]),.b(fsu[191]),.cin(fca[182]),.sum(fsu[426]),.carry(fca[426]));
FA FA427 (.a(fsu[192]),.b(fca[183]),.cin(pp[4][30]),.sum(fsu[427]),.carry(fca[427]));
FA FA428 (.a(fca[184]),.b(fsu[193]),.cin(fca[185]),.sum(fsu[428]),.carry(fca[428]));
FA FA429 (.a(fsu[194]),.b(fca[186]),.cin(fsu[195]),.sum(fsu[429]),.carry(fca[429]));
FA FA430 (.a(fca[187]),.b(fsu[196]),.cin(fca[188]),.sum(fsu[430]),.carry(fca[430]));
FA FA431 (.a(fsu[197]),.b(fca[189]),.cin(fsu[198]),.sum(fsu[431]),.carry(fca[431]));
FA FA432 (.a(fca[190]),.b(fsu[199]),.cin(fca[191]),.sum(fsu[432]),.carry(fca[432]));
FA FA433 (.a(fsu[200]),.b(fca[192]),.cin(pp[5][30]),.sum(fsu[433]),.carry(fca[433]));
FA FA434 (.a(hca[12]),.b(fsu[201]),.cin(fca[193]),.sum(fsu[434]),.carry(fca[434]));
FA FA435 (.a(fsu[202]),.b(fca[194]),.cin(fsu[203]),.sum(fsu[435]),.carry(fca[435]));
FA FA436 (.a(fca[195]),.b(fsu[204]),.cin(fca[196]),.sum(fsu[436]),.carry(fca[436]));
FA FA437 (.a(fsu[205]),.b(fca[197]),.cin(fsu[206]),.sum(fsu[437]),.carry(fca[437]));
FA FA438 (.a(fca[198]),.b(fsu[207]),.cin(fca[199]),.sum(fsu[438]),.carry(fca[438]));
FA FA439 (.a(fsu[208]),.b(fca[200]),.cin(pp[6][30]),.sum(fsu[439]),.carry(fca[439]));
HA HA31 (.a(fsu[209]),.b(fca[201]),.sum_h(hsu[31]),.carry_h(hca[31]));
FA FA440 (.a(fsu[210]),.b(fca[202]),.cin(fsu[211]),.sum(fsu[440]),.carry(fca[440]));
FA FA441 (.a(fca[203]),.b(fsu[212]),.cin(fca[204]),.sum(fsu[441]),.carry(fca[441]));
FA FA442 (.a(fsu[213]),.b(fca[205]),.cin(fsu[214]),.sum(fsu[442]),.carry(fca[442]));
FA FA443 (.a(fca[206]),.b(fsu[215]),.cin(fca[207]),.sum(fsu[443]),.carry(fca[443]));
FA FA444 (.a(fsu[216]),.b(fca[208]),.cin(pp[7][30]),.sum(fsu[444]),.carry(fca[444]));
HA HA32 (.a(hsu[13]),.b(fca[209]),.sum_h(hsu[32]),.carry_h(hca[32]));
FA FA445 (.a(fsu[217]),.b(fca[210]),.cin(fsu[218]),.sum(fsu[445]),.carry(fca[445]));
FA FA446 (.a(fca[211]),.b(fsu[219]),.cin(fca[212]),.sum(fsu[446]),.carry(fca[446]));
FA FA447 (.a(fsu[220]),.b(fca[213]),.cin(fsu[221]),.sum(fsu[447]),.carry(fca[447]));
FA FA448 (.a(fca[214]),.b(fsu[222]),.cin(fca[215]),.sum(fsu[448]),.carry(fca[448]));
FA FA449 (.a(fsu[223]),.b(fca[216]),.cin(pp[8][30]),.sum(fsu[449]),.carry(fca[449]));
HA HA33 (.a(pp[31][8]),.b(hca[13]),.sum_h(hsu[33]),.carry_h(hca[33]));
FA FA450 (.a(fsu[224]),.b(fca[217]),.cin(fsu[225]),.sum(fsu[450]),.carry(fca[450]));
FA FA451 (.a(fca[218]),.b(fsu[226]),.cin(fca[219]),.sum(fsu[451]),.carry(fca[451]));
FA FA452 (.a(fsu[227]),.b(fca[220]),.cin(fsu[228]),.sum(fsu[452]),.carry(fca[452]));
FA FA453 (.a(fca[221]),.b(fsu[229]),.cin(fca[222]),.sum(fsu[453]),.carry(fca[453]));
FA FA454 (.a(fsu[230]),.b(fca[223]),.cin(pp[9][30]),.sum(fsu[454]),.carry(fca[454]));
FA FA455 (.a(fsu[231]),.b(fca[224]),.cin(fsu[232]),.sum(fsu[455]),.carry(fca[455]));
FA FA456 (.a(fca[225]),.b(fsu[233]),.cin(fca[226]),.sum(fsu[456]),.carry(fca[456]));
FA FA457 (.a(fsu[234]),.b(fca[227]),.cin(fsu[235]),.sum(fsu[457]),.carry(fca[457]));
FA FA458 (.a(fca[228]),.b(fsu[236]),.cin(fca[229]),.sum(fsu[458]),.carry(fca[458]));
FA FA459 (.a(fsu[237]),.b(fca[230]),.cin(pp[10][30]),.sum(fsu[459]),.carry(fca[459]));
FA FA460 (.a(hsu[14]),.b(fca[231]),.cin(fsu[238]),.sum(fsu[460]),.carry(fca[460]));
FA FA461 (.a(fca[232]),.b(fsu[239]),.cin(fca[233]),.sum(fsu[461]),.carry(fca[461]));
FA FA462 (.a(fsu[240]),.b(fca[234]),.cin(fsu[241]),.sum(fsu[462]),.carry(fca[462]));
FA FA463 (.a(fca[235]),.b(fsu[242]),.cin(fca[236]),.sum(fsu[463]),.carry(fca[463]));
FA FA464 (.a(fsu[243]),.b(fca[237]),.cin(pp[11][30]),.sum(fsu[464]),.carry(fca[464]));
FA FA465 (.a(pp[31][11]),.b(hca[14]),.cin(fsu[244]),.sum(fsu[465]),.carry(fca[465]));
FA FA466 (.a(fca[238]),.b(fsu[245]),.cin(fca[239]),.sum(fsu[466]),.carry(fca[466]));
FA FA467 (.a(fsu[246]),.b(fca[240]),.cin(fsu[247]),.sum(fsu[467]),.carry(fca[467]));
FA FA468 (.a(fca[241]),.b(fsu[248]),.cin(fca[242]),.sum(fsu[468]),.carry(fca[468]));
FA FA469 (.a(fsu[249]),.b(fca[243]),.cin(pp[12][30]),.sum(fsu[469]),.carry(fca[469]));
FA FA470 (.a(fca[244]),.b(fsu[251]),.cin(fca[245]),.sum(fsu[470]),.carry(fca[470]));
FA FA471 (.a(fsu[252]),.b(fca[246]),.cin(fsu[253]),.sum(fsu[471]),.carry(fca[471]));
FA FA472 (.a(fca[247]),.b(fsu[254]),.cin(fca[248]),.sum(fsu[472]),.carry(fca[472]));
FA FA473 (.a(fsu[255]),.b(fca[249]),.cin(pp[13][30]),.sum(fsu[473]),.carry(fca[473]));
FA FA474 (.a(fca[250]),.b(fsu[256]),.cin(fca[251]),.sum(fsu[474]),.carry(fca[474]));
FA FA475 (.a(fsu[257]),.b(fca[252]),.cin(fsu[258]),.sum(fsu[475]),.carry(fca[475]));
FA FA476 (.a(fca[253]),.b(fsu[259]),.cin(fca[254]),.sum(fsu[476]),.carry(fca[476]));
FA FA477 (.a(fsu[260]),.b(fca[255]),.cin(pp[14][30]),.sum(fsu[477]),.carry(fca[477]));
FA FA478 (.a(hca[15]),.b(fsu[261]),.cin(fca[256]),.sum(fsu[478]),.carry(fca[478]));
FA FA479 (.a(fsu[262]),.b(fca[257]),.cin(fsu[263]),.sum(fsu[479]),.carry(fca[479]));
FA FA480 (.a(fca[258]),.b(fsu[264]),.cin(fca[259]),.sum(fsu[480]),.carry(fca[480]));
FA FA481 (.a(fsu[265]),.b(fca[260]),.cin(pp[15][30]),.sum(fsu[481]),.carry(fca[481]));
HA HA34 (.a(fsu[266]),.b(fca[261]),.sum_h(hsu[34]),.carry_h(hca[34]));
FA FA482 (.a(fsu[267]),.b(fca[262]),.cin(fsu[268]),.sum(fsu[482]),.carry(fca[482]));
FA FA483 (.a(fca[263]),.b(fsu[269]),.cin(fca[264]),.sum(fsu[483]),.carry(fca[483]));
FA FA484 (.a(fsu[270]),.b(fca[265]),.cin(pp[16][30]),.sum(fsu[484]),.carry(fca[484]));
HA HA35 (.a(hsu[16]),.b(fca[266]),.sum_h(hsu[35]),.carry_h(hca[35]));
FA FA485 (.a(fsu[271]),.b(fca[267]),.cin(fsu[272]),.sum(fsu[485]),.carry(fca[485]));
FA FA486 (.a(fca[268]),.b(fsu[273]),.cin(fca[269]),.sum(fsu[486]),.carry(fca[486]));
FA FA487 (.a(fsu[274]),.b(fca[270]),.cin(pp[17][30]),.sum(fsu[487]),.carry(fca[487]));
HA HA36 (.a(pp[31][17]),.b(hca[16]),.sum_h(hsu[36]),.carry_h(hca[36]));
FA FA488 (.a(fsu[275]),.b(fca[271]),.cin(fsu[276]),.sum(fsu[488]),.carry(fca[488]));
FA FA489 (.a(fca[272]),.b(fsu[277]),.cin(fca[273]),.sum(fsu[489]),.carry(fca[489]));
FA FA490 (.a(fsu[278]),.b(fca[274]),.cin(pp[18][30]),.sum(fsu[490]),.carry(fca[490]));
FA FA491 (.a(fsu[279]),.b(fca[275]),.cin(fsu[280]),.sum(fsu[491]),.carry(fca[491]));
FA FA492 (.a(fca[276]),.b(fsu[281]),.cin(fca[277]),.sum(fsu[492]),.carry(fca[492]));
FA FA493 (.a(fsu[282]),.b(fca[278]),.cin(pp[19][30]),.sum(fsu[493]),.carry(fca[493]));
FA FA494 (.a(hsu[17]),.b(fca[279]),.cin(fsu[283]),.sum(fsu[494]),.carry(fca[494]));
FA FA495 (.a(fca[280]),.b(fsu[284]),.cin(fca[281]),.sum(fsu[495]),.carry(fca[495]));
FA FA496 (.a(fsu[285]),.b(fca[282]),.cin(pp[20][30]),.sum(fsu[496]),.carry(fca[496]));
FA FA497 (.a(pp[31][20]),.b(hca[17]),.cin(fsu[286]),.sum(fsu[497]),.carry(fca[497]));
FA FA498 (.a(fca[283]),.b(fsu[287]),.cin(fca[284]),.sum(fsu[498]),.carry(fca[498]));
FA FA499 (.a(fsu[288]),.b(fca[285]),.cin(pp[21][30]),.sum(fsu[499]),.carry(fca[499]));
FA FA500 (.a(fca[286]),.b(fsu[290]),.cin(fca[287]),.sum(fsu[500]),.carry(fca[500]));
FA FA501 (.a(fsu[291]),.b(fca[288]),.cin(pp[22][30]),.sum(fsu[501]),.carry(fca[501]));
FA FA502 (.a(fca[289]),.b(fsu[292]),.cin(fca[290]),.sum(fsu[502]),.carry(fca[502]));
FA FA503 (.a(fsu[293]),.b(fca[291]),.cin(pp[23][30]),.sum(fsu[503]),.carry(fca[503]));
FA FA504 (.a(hca[18]),.b(fsu[294]),.cin(fca[292]),.sum(fsu[504]),.carry(fca[504]));
FA FA505 (.a(fsu[295]),.b(fca[293]),.cin(pp[24][30]),.sum(fsu[505]),.carry(fca[505]));
HA HA37 (.a(fsu[296]),.b(fca[294]),.sum_h(hsu[37]),.carry_h(hca[37]));
FA FA506 (.a(fsu[297]),.b(fca[295]),.cin(pp[25][30]),.sum(fsu[506]),.carry(fca[506]));
HA HA38 (.a(hsu[19]),.b(fca[296]),.sum_h(hsu[38]),.carry_h(hca[38]));
FA FA507 (.a(fsu[298]),.b(fca[297]),.cin(pp[26][30]),.sum(fsu[507]),.carry(fca[507]));
HA HA39 (.a(pp[31][26]),.b(hca[19]),.sum_h(hsu[39]),.carry_h(hca[39]));
FA FA508 (.a(fsu[299]),.b(fca[298]),.cin(pp[27][30]),.sum(fsu[508]),.carry(fca[508]));
FA FA509 (.a(fsu[300]),.b(fca[299]),.cin(pp[28][30]),.sum(fsu[509]),.carry(fca[509]));
FA FA510 (.a(hsu[20]),.b(fca[300]),.cin(pp[29][30]),.sum(fsu[510]),.carry(fca[510]));
FA FA511 (.a(pp[31][29]),.b(hca[20]),.cin(pp[30][30]),.sum(fsu[511]),.carry(fca[511]));
//3rd stage
HA HA40 (.a(fsu[301]),.b(hca[21]),.sum_h(z[3]),.carry_h(hca[40]));
HA HA41 (.a(fsu[302]),.b(fca[301]),.sum_h(hsu[41]),.carry_h(hca[41]));
FA FA512 (.a(fsu[303]),.b(fca[302]),.cin(hca[2]),.sum(fsu[512]),.carry(fca[512]));
FA FA513 (.a(fsu[304]),.b(fca[303]),.cin(hsu[22]),.sum(fsu[513]),.carry(fca[513]));
FA FA514 (.a(fsu[305]),.b(fca[304]),.cin(hsu[23]),.sum(fsu[514]),.carry(fca[514]));
FA FA515 (.a(fsu[306]),.b(fca[305]),.cin(fsu[307]),.sum(fsu[515]),.carry(fca[515]));
FA FA516 (.a(fsu[308]),.b(fca[306]),.cin(fsu[309]),.sum(fsu[516]),.carry(fca[516]));
HA HA42 (.a(fca[307]),.b(pp[0][9]),.sum_h(hsu[42]),.carry_h(hca[42]));
FA FA517 (.a(fsu[310]),.b(fca[308]),.cin(fsu[311]),.sum(fsu[517]),.carry(fca[517]));
HA HA43 (.a(fca[309]),.b(hsu[4]),.sum_h(hsu[43]),.carry_h(hca[43]));
FA FA518 (.a(fsu[312]),.b(fca[310]),.cin(fsu[313]),.sum(fsu[518]),.carry(fca[518]));
HA HA44 (.a(fca[311]),.b(hsu[24]),.sum_h(hsu[44]),.carry_h(hca[44]));
FA FA519 (.a(fsu[314]),.b(fca[312]),.cin(fsu[315]),.sum(fsu[519]),.carry(fca[519]));
FA FA520 (.a(fca[313]),.b(fsu[316]),.cin(hca[24]),.sum(fsu[520]),.carry(fca[520]));
FA FA521 (.a(fsu[317]),.b(fca[314]),.cin(fsu[318]),.sum(fsu[521]),.carry(fca[521]));
FA FA522 (.a(fca[315]),.b(fsu[319]),.cin(fca[316]),.sum(fsu[522]),.carry(fca[522]));
FA FA523 (.a(fsu[320]),.b(fca[317]),.cin(fsu[321]),.sum(fsu[523]),.carry(fca[523]));
FA FA524 (.a(fca[318]),.b(fsu[322]),.cin(fca[319]),.sum(fsu[524]),.carry(fca[524]));
FA FA525 (.a(fsu[323]),.b(fca[320]),.cin(fsu[324]),.sum(fsu[525]),.carry(fca[525]));
FA FA526 (.a(fca[321]),.b(fsu[325]),.cin(fca[322]),.sum(fsu[526]),.carry(fca[526]));
FA FA527 (.a(fsu[326]),.b(fca[323]),.cin(fsu[327]),.sum(fsu[527]),.carry(fca[527]));
FA FA528 (.a(fca[324]),.b(fsu[328]),.cin(fca[325]),.sum(fsu[528]),.carry(fca[528]));
HA HA45 (.a(hsu[26]),.b(hca[25]),.sum_h(hsu[45]),.carry_h(hca[45]));
FA FA529 (.a(fsu[329]),.b(fca[326]),.cin(fsu[330]),.sum(fsu[529]),.carry(fca[529]));
FA FA530 (.a(fca[327]),.b(fsu[331]),.cin(fca[328]),.sum(fsu[530]),.carry(fca[530]));
HA HA46 (.a(fsu[332]),.b(hca[26]),.sum_h(hsu[46]),.carry_h(hca[46]));
FA FA531 (.a(fsu[333]),.b(fca[329]),.cin(fsu[334]),.sum(fsu[531]),.carry(fca[531]));
FA FA532 (.a(fca[330]),.b(fsu[335]),.cin(fca[331]),.sum(fsu[532]),.carry(fca[532]));
FA FA533 (.a(fsu[336]),.b(fca[332]),.cin(pp[0][18]),.sum(fsu[533]),.carry(fca[533]));
FA FA534 (.a(fsu[337]),.b(fca[333]),.cin(fsu[338]),.sum(fsu[534]),.carry(fca[534]));
FA FA535 (.a(fca[334]),.b(fsu[339]),.cin(fca[335]),.sum(fsu[535]),.carry(fca[535]));
FA FA536 (.a(fsu[340]),.b(fca[336]),.cin(hsu[7]),.sum(fsu[536]),.carry(fca[536]));
FA FA537 (.a(fsu[341]),.b(fca[337]),.cin(fsu[342]),.sum(fsu[537]),.carry(fca[537]));
FA FA538 (.a(fca[338]),.b(fsu[343]),.cin(fca[339]),.sum(fsu[538]),.carry(fca[538]));
FA FA539 (.a(fsu[344]),.b(fca[340]),.cin(hsu[27]),.sum(fsu[539]),.carry(fca[539]));
FA FA540 (.a(fsu[345]),.b(fca[341]),.cin(fsu[346]),.sum(fsu[540]),.carry(fca[540]));
FA FA541 (.a(fca[342]),.b(fsu[347]),.cin(fca[343]),.sum(fsu[541]),.carry(fca[541]));
FA FA542 (.a(fsu[348]),.b(fca[344]),.cin(fsu[349]),.sum(fsu[542]),.carry(fca[542]));
FA FA543 (.a(fsu[350]),.b(fca[345]),.cin(fsu[351]),.sum(fsu[543]),.carry(fca[543]));
FA FA544 (.a(fca[346]),.b(fsu[352]),.cin(fca[347]),.sum(fsu[544]),.carry(fca[544]));
FA FA545 (.a(fsu[353]),.b(fca[348]),.cin(fsu[354]),.sum(fsu[545]),.carry(fca[545]));
FA FA546 (.a(fsu[355]),.b(fca[350]),.cin(fsu[356]),.sum(fsu[546]),.carry(fca[546]));
FA FA547 (.a(fca[351]),.b(fsu[357]),.cin(fca[352]),.sum(fsu[547]),.carry(fca[547]));
FA FA548 (.a(fsu[358]),.b(fca[353]),.cin(fsu[359]),.sum(fsu[548]),.carry(fca[548]));
HA HA47 (.a(fca[354]),.b(hca[8]),.sum_h(hsu[47]),.carry_h(hca[47]));
FA FA549 (.a(fsu[360]),.b(fca[355]),.cin(fsu[361]),.sum(fsu[549]),.carry(fca[549]));
FA FA550 (.a(fca[356]),.b(fsu[362]),.cin(fca[357]),.sum(fsu[550]),.carry(fca[550]));
FA FA551 (.a(fsu[363]),.b(fca[358]),.cin(fsu[364]),.sum(fsu[551]),.carry(fca[551]));
HA HA48 (.a(fca[359]),.b(hsu[28]),.sum_h(hsu[48]),.carry_h(hca[48]));
FA FA552 (.a(fsu[365]),.b(fca[360]),.cin(fsu[366]),.sum(fsu[552]),.carry(fca[552]));
FA FA553 (.a(fca[361]),.b(fsu[367]),.cin(fca[362]),.sum(fsu[553]),.carry(fca[553]));
FA FA554 (.a(fsu[368]),.b(fca[363]),.cin(fsu[369]),.sum(fsu[554]),.carry(fca[554]));
FA FA555 (.a(fca[364]),.b(hsu[29]),.cin(hca[28]),.sum(fsu[555]),.carry(fca[555]));
FA FA556 (.a(fsu[370]),.b(fca[365]),.cin(fsu[371]),.sum(fsu[556]),.carry(fca[556]));
FA FA557 (.a(fca[366]),.b(fsu[372]),.cin(fca[367]),.sum(fsu[557]),.carry(fca[557]));
FA FA558 (.a(fsu[373]),.b(fca[368]),.cin(fsu[374]),.sum(fsu[558]),.carry(fca[558]));
FA FA559 (.a(fca[369]),.b(fsu[375]),.cin(hca[29]),.sum(fsu[559]),.carry(fca[559]));
FA FA560 (.a(fsu[376]),.b(fca[370]),.cin(fsu[377]),.sum(fsu[560]),.carry(fca[560]));
FA FA561 (.a(fca[371]),.b(fsu[378]),.cin(fca[372]),.sum(fsu[561]),.carry(fca[561]));
FA FA562 (.a(fsu[379]),.b(fca[373]),.cin(fsu[380]),.sum(fsu[562]),.carry(fca[562]));
FA FA563 (.a(fca[374]),.b(fsu[381]),.cin(fca[375]),.sum(fsu[563]),.carry(fca[563]));
FA FA564 (.a(fsu[382]),.b(fca[376]),.cin(fsu[383]),.sum(fsu[564]),.carry(fca[564]));
FA FA565 (.a(fca[377]),.b(fsu[384]),.cin(fca[378]),.sum(fsu[565]),.carry(fca[565]));
FA FA566 (.a(fsu[385]),.b(fca[379]),.cin(fsu[386]),.sum(fsu[566]),.carry(fca[566]));
FA FA567 (.a(fca[380]),.b(fsu[387]),.cin(fca[381]),.sum(fsu[567]),.carry(fca[567]));
FA FA568 (.a(fsu[388]),.b(fca[382]),.cin(fsu[389]),.sum(fsu[568]),.carry(fca[568]));
FA FA569 (.a(fca[383]),.b(fsu[390]),.cin(fca[384]),.sum(fsu[569]),.carry(fca[569]));
FA FA570 (.a(fsu[391]),.b(fca[385]),.cin(fsu[392]),.sum(fsu[570]),.carry(fca[570]));
FA FA571 (.a(fca[386]),.b(fsu[393]),.cin(fca[387]),.sum(fsu[571]),.carry(fca[571]));
FA FA572 (.a(fsu[394]),.b(fca[388]),.cin(fsu[395]),.sum(fsu[572]),.carry(fca[572]));
FA FA573 (.a(fca[389]),.b(fsu[396]),.cin(fca[390]),.sum(fsu[573]),.carry(fca[573]));
FA FA574 (.a(fsu[397]),.b(fca[391]),.cin(fsu[398]),.sum(fsu[574]),.carry(fca[574]));
FA FA575 (.a(fca[392]),.b(fsu[399]),.cin(fca[393]),.sum(fsu[575]),.carry(fca[575]));
HA HA49 (.a(fsu[400]),.b(hca[30]),.sum_h(hsu[49]),.carry_h(hca[49]));
FA FA576 (.a(fsu[401]),.b(fca[394]),.cin(fsu[402]),.sum(fsu[576]),.carry(fca[576]));
FA FA577 (.a(fca[395]),.b(fsu[403]),.cin(fca[396]),.sum(fsu[577]),.carry(fca[577]));
FA FA578 (.a(fsu[404]),.b(fca[397]),.cin(fsu[405]),.sum(fsu[578]),.carry(fca[578]));
FA FA579 (.a(fca[398]),.b(fsu[406]),.cin(fca[399]),.sum(fsu[579]),.carry(fca[579]));
FA FA580 (.a(fsu[407]),.b(fca[400]),.cin(pp[0][31]),.sum(fsu[580]),.carry(fca[580]));
FA FA581 (.a(fsu[408]),.b(fca[401]),.cin(fsu[409]),.sum(fsu[581]),.carry(fca[581]));
FA FA582 (.a(fca[402]),.b(fsu[410]),.cin(fca[403]),.sum(fsu[582]),.carry(fca[582]));
FA FA583 (.a(fsu[411]),.b(fca[404]),.cin(fsu[412]),.sum(fsu[583]),.carry(fca[583]));
FA FA584 (.a(fca[405]),.b(fsu[413]),.cin(fca[406]),.sum(fsu[584]),.carry(fca[584]));
FA FA585 (.a(fsu[414]),.b(fca[407]),.cin(pp[1][31]),.sum(fsu[585]),.carry(fca[585]));
FA FA586 (.a(fsu[415]),.b(fca[408]),.cin(fsu[416]),.sum(fsu[586]),.carry(fca[586]));
FA FA587 (.a(fca[409]),.b(fsu[417]),.cin(fca[410]),.sum(fsu[587]),.carry(fca[587]));
FA FA588 (.a(fsu[418]),.b(fca[411]),.cin(fsu[419]),.sum(fsu[588]),.carry(fca[588]));
FA FA589 (.a(fca[412]),.b(fsu[420]),.cin(fca[413]),.sum(fsu[589]),.carry(fca[589]));
FA FA590 (.a(fsu[421]),.b(fca[414]),.cin(pp[2][31]),.sum(fsu[590]),.carry(fca[590]));
FA FA591 (.a(fsu[184]),.b(fca[415]),.cin(fsu[422]),.sum(fsu[591]),.carry(fca[591]));
FA FA592 (.a(fca[416]),.b(fsu[423]),.cin(fca[417]),.sum(fsu[592]),.carry(fca[592]));
FA FA593 (.a(fsu[424]),.b(fca[418]),.cin(fsu[425]),.sum(fsu[593]),.carry(fca[593]));
FA FA594 (.a(fca[419]),.b(fsu[426]),.cin(fca[420]),.sum(fsu[594]),.carry(fca[594]));
FA FA595 (.a(fsu[427]),.b(fca[421]),.cin(pp[3][31]),.sum(fsu[595]),.carry(fca[595]));
HA HA50 (.a(hsu[12]),.b(fsu[428]),.sum_h(hsu[50]),.carry_h(hca[50]));
FA FA596 (.a(fca[422]),.b(fsu[429]),.cin(fca[423]),.sum(fsu[596]),.carry(fca[596]));
FA FA597 (.a(fsu[430]),.b(fca[424]),.cin(fsu[431]),.sum(fsu[597]),.carry(fca[597]));
FA FA598 (.a(fca[425]),.b(fsu[432]),.cin(fca[426]),.sum(fsu[598]),.carry(fca[598]));
FA FA599 (.a(fsu[433]),.b(fca[427]),.cin(pp[4][31]),.sum(fsu[599]),.carry(fca[599]));
HA HA51 (.a(pp[31][5]),.b(fsu[434]),.sum_h(hsu[51]),.carry_h(hca[51]));
FA FA600 (.a(fca[428]),.b(fsu[435]),.cin(fca[429]),.sum(fsu[600]),.carry(fca[600]));
FA FA601 (.a(fsu[436]),.b(fca[430]),.cin(fsu[437]),.sum(fsu[601]),.carry(fca[601]));
FA FA602 (.a(fca[431]),.b(fsu[438]),.cin(fca[432]),.sum(fsu[602]),.carry(fca[602]));
FA FA603 (.a(fsu[439]),.b(fca[433]),.cin(pp[5][31]),.sum(fsu[603]),.carry(fca[603]));
FA FA604 (.a(fca[434]),.b(fsu[440]),.cin(fca[435]),.sum(fsu[604]),.carry(fca[604]));
FA FA605 (.a(fsu[441]),.b(fca[436]),.cin(fsu[442]),.sum(fsu[605]),.carry(fca[605]));
FA FA606 (.a(fca[437]),.b(fsu[443]),.cin(fca[438]),.sum(fsu[606]),.carry(fca[606]));
FA FA607 (.a(fsu[444]),.b(fca[439]),.cin(pp[6][31]),.sum(fsu[607]),.carry(fca[607]));
FA FA608 (.a(hca[31]),.b(fsu[445]),.cin(fca[440]),.sum(fsu[608]),.carry(fca[608]));
FA FA609 (.a(fsu[446]),.b(fca[441]),.cin(fsu[447]),.sum(fsu[609]),.carry(fca[609]));
FA FA610 (.a(fca[442]),.b(fsu[448]),.cin(fca[443]),.sum(fsu[610]),.carry(fca[610]));
FA FA611 (.a(fsu[449]),.b(fca[444]),.cin(pp[7][31]),.sum(fsu[611]),.carry(fca[611]));
FA FA612 (.a(hca[32]),.b(fsu[450]),.cin(fca[445]),.sum(fsu[612]),.carry(fca[612]));
FA FA613 (.a(fsu[451]),.b(fca[446]),.cin(fsu[452]),.sum(fsu[613]),.carry(fca[613]));
FA FA614 (.a(fca[447]),.b(fsu[453]),.cin(fca[448]),.sum(fsu[614]),.carry(fca[614]));
FA FA615 (.a(fsu[454]),.b(fca[449]),.cin(pp[8][31]),.sum(fsu[615]),.carry(fca[615]));
FA FA616 (.a(hca[33]),.b(fsu[455]),.cin(fca[450]),.sum(fsu[616]),.carry(fca[616]));
FA FA617 (.a(fsu[456]),.b(fca[451]),.cin(fsu[457]),.sum(fsu[617]),.carry(fca[617]));
FA FA618 (.a(fca[452]),.b(fsu[458]),.cin(fca[453]),.sum(fsu[618]),.carry(fca[618]));
FA FA619 (.a(fsu[459]),.b(fca[454]),.cin(pp[9][31]),.sum(fsu[619]),.carry(fca[619]));
HA HA52 (.a(fsu[460]),.b(fca[455]),.sum_h(hsu[52]),.carry_h(hca[52]));
FA FA620 (.a(fsu[461]),.b(fca[456]),.cin(fsu[462]),.sum(fsu[620]),.carry(fca[620]));
FA FA621 (.a(fca[457]),.b(fsu[463]),.cin(fca[458]),.sum(fsu[621]),.carry(fca[621]));
FA FA622 (.a(fsu[464]),.b(fca[459]),.cin(pp[10][31]),.sum(fsu[622]),.carry(fca[622]));
HA HA53 (.a(fsu[465]),.b(fca[460]),.sum_h(hsu[53]),.carry_h(hca[53]));
FA FA623 (.a(fsu[466]),.b(fca[461]),.cin(fsu[467]),.sum(fsu[623]),.carry(fca[623]));
FA FA624 (.a(fca[462]),.b(fsu[468]),.cin(fca[463]),.sum(fsu[624]),.carry(fca[624]));
FA FA625 (.a(fsu[469]),.b(fca[464]),.cin(pp[11][31]),.sum(fsu[625]),.carry(fca[625]));
HA HA54 (.a(fsu[250]),.b(fca[465]),.sum_h(hsu[54]),.carry_h(hca[54]));
FA FA626 (.a(fsu[470]),.b(fca[466]),.cin(fsu[471]),.sum(fsu[626]),.carry(fca[626]));
FA FA627 (.a(fca[467]),.b(fsu[472]),.cin(fca[468]),.sum(fsu[627]),.carry(fca[627]));
FA FA628 (.a(fsu[473]),.b(fca[469]),.cin(pp[12][31]),.sum(fsu[628]),.carry(fca[628]));
FA FA629 (.a(fsu[474]),.b(fca[470]),.cin(fsu[475]),.sum(fsu[629]),.carry(fca[629]));
FA FA630 (.a(fca[471]),.b(fsu[476]),.cin(fca[472]),.sum(fsu[630]),.carry(fca[630]));
FA FA631 (.a(fsu[477]),.b(fca[473]),.cin(pp[13][31]),.sum(fsu[631]),.carry(fca[631]));
FA FA632 (.a(fsu[478]),.b(fca[474]),.cin(fsu[479]),.sum(fsu[632]),.carry(fca[632]));
FA FA633 (.a(fca[475]),.b(fsu[480]),.cin(fca[476]),.sum(fsu[633]),.carry(fca[633]));
FA FA634 (.a(fsu[481]),.b(fca[477]),.cin(pp[14][31]),.sum(fsu[634]),.carry(fca[634]));
FA FA635 (.a(hsu[34]),.b(fca[478]),.cin(fsu[482]),.sum(fsu[635]),.carry(fca[635]));
FA FA636 (.a(fca[479]),.b(fsu[483]),.cin(fca[480]),.sum(fsu[636]),.carry(fca[636]));
FA FA637 (.a(fsu[484]),.b(fca[481]),.cin(pp[15][31]),.sum(fsu[637]),.carry(fca[637]));
FA FA638 (.a(hsu[35]),.b(hca[34]),.cin(fsu[485]),.sum(fsu[638]),.carry(fca[638]));
FA FA639 (.a(fca[482]),.b(fsu[486]),.cin(fca[483]),.sum(fsu[639]),.carry(fca[639]));
FA FA640 (.a(fsu[487]),.b(fca[484]),.cin(pp[16][31]),.sum(fsu[640]),.carry(fca[640]));
FA FA641 (.a(hsu[36]),.b(hca[35]),.cin(fsu[488]),.sum(fsu[641]),.carry(fca[641]));
FA FA642 (.a(fca[485]),.b(fsu[489]),.cin(fca[486]),.sum(fsu[642]),.carry(fca[642]));
FA FA643 (.a(fsu[490]),.b(fca[487]),.cin(pp[17][31]),.sum(fsu[643]),.carry(fca[643]));
HA HA55 (.a(hca[36]),.b(fsu[491]),.sum_h(hsu[55]),.carry_h(hca[55]));
FA FA644 (.a(fca[488]),.b(fsu[492]),.cin(fca[489]),.sum(fsu[644]),.carry(fca[644]));
FA FA645 (.a(fsu[493]),.b(fca[490]),.cin(pp[18][31]),.sum(fsu[645]),.carry(fca[645]));
FA FA646 (.a(fca[491]),.b(fsu[495]),.cin(fca[492]),.sum(fsu[646]),.carry(fca[646]));
FA FA647 (.a(fsu[496]),.b(fca[493]),.cin(pp[19][31]),.sum(fsu[647]),.carry(fca[647]));
FA FA648 (.a(fca[494]),.b(fsu[498]),.cin(fca[495]),.sum(fsu[648]),.carry(fca[648]));
FA FA649 (.a(fsu[499]),.b(fca[496]),.cin(pp[20][31]),.sum(fsu[649]),.carry(fca[649]));
FA FA650 (.a(fca[497]),.b(fsu[500]),.cin(fca[498]),.sum(fsu[650]),.carry(fca[650]));
FA FA651 (.a(fsu[501]),.b(fca[499]),.cin(pp[21][31]),.sum(fsu[651]),.carry(fca[651]));
FA FA652 (.a(hsu[18]),.b(fsu[502]),.cin(fca[500]),.sum(fsu[652]),.carry(fca[652]));
FA FA653 (.a(fsu[503]),.b(fca[501]),.cin(pp[22][31]),.sum(fsu[653]),.carry(fca[653]));
FA FA654 (.a(pp[31][23]),.b(fsu[504]),.cin(fca[502]),.sum(fsu[654]),.carry(fca[654]));
FA FA655 (.a(fsu[505]),.b(fca[503]),.cin(pp[23][31]),.sum(fsu[655]),.carry(fca[655]));
HA HA56 (.a(hsu[37]),.b(fca[504]),.sum_h(hsu[56]),.carry_h(hca[56]));
FA FA656 (.a(fsu[506]),.b(fca[505]),.cin(pp[24][31]),.sum(fsu[656]),.carry(fca[656]));
HA HA57 (.a(hsu[38]),.b(hca[37]),.sum_h(hsu[57]),.carry_h(hca[57]));
FA FA657 (.a(fsu[507]),.b(fca[506]),.cin(pp[25][31]),.sum(fsu[657]),.carry(fca[657]));
HA HA58 (.a(hsu[39]),.b(hca[38]),.sum_h(hsu[58]),.carry_h(hca[58]));
FA FA658 (.a(fsu[508]),.b(fca[507]),.cin(pp[26][31]),.sum(fsu[658]),.carry(fca[658]));
FA FA659 (.a(fsu[509]),.b(fca[508]),.cin(pp[27][31]),.sum(fsu[659]),.carry(fca[659]));
FA FA660 (.a(fsu[510]),.b(fca[509]),.cin(pp[28][31]),.sum(fsu[660]),.carry(fca[660]));
FA FA661 (.a(fsu[511]),.b(fca[510]),.cin(pp[29][31]),.sum(fsu[661]),.carry(fca[661]));
FA FA662 (.a(pp[31][30]),.b(fca[511]),.cin(pp[30][31]),.sum(fsu[662]),.carry(fca[662]));
//4th stage
HA HA59 (.a(hsu[41]),.b(hca[40]),.sum_h(z[4]),.carry_h(hca[59]));
HA HA60 (.a(fsu[512]),.b(hca[41]),.sum_h(hsu[60]),.carry_h(hca[60]));
HA HA61 (.a(fsu[513]),.b(fca[512]),.sum_h(hsu[61]),.carry_h(hca[61]));
FA FA663 (.a(fsu[514]),.b(fca[513]),.cin(hca[22]),.sum(fsu[663]),.carry(fca[663]));
FA FA664 (.a(fsu[515]),.b(fca[514]),.cin(hca[23]),.sum(fsu[664]),.carry(fca[664]));
FA FA665 (.a(fsu[516]),.b(fca[515]),.cin(hsu[42]),.sum(fsu[665]),.carry(fca[665]));
FA FA666 (.a(fsu[517]),.b(fca[516]),.cin(hsu[43]),.sum(fsu[666]),.carry(fca[666]));
FA FA667 (.a(fsu[518]),.b(fca[517]),.cin(hsu[44]),.sum(fsu[667]),.carry(fca[667]));
FA FA668 (.a(fsu[519]),.b(fca[518]),.cin(fsu[520]),.sum(fsu[668]),.carry(fca[668]));
FA FA669 (.a(fsu[521]),.b(fca[519]),.cin(fsu[522]),.sum(fsu[669]),.carry(fca[669]));
FA FA670 (.a(fsu[523]),.b(fca[521]),.cin(fsu[524]),.sum(fsu[670]),.carry(fca[670]));
HA HA62 (.a(fca[522]),.b(hca[5]),.sum_h(hsu[62]),.carry_h(hca[62]));
FA FA671 (.a(fsu[525]),.b(fca[523]),.cin(fsu[526]),.sum(fsu[671]),.carry(fca[671]));
HA HA63 (.a(fca[524]),.b(hsu[25]),.sum_h(hsu[63]),.carry_h(hca[63]));
FA FA672 (.a(fsu[527]),.b(fca[525]),.cin(fsu[528]),.sum(fsu[672]),.carry(fca[672]));
HA HA64 (.a(fca[526]),.b(hsu[45]),.sum_h(hsu[64]),.carry_h(hca[64]));
FA FA673 (.a(fsu[529]),.b(fca[527]),.cin(fsu[530]),.sum(fsu[673]),.carry(fca[673]));
FA FA674 (.a(fca[528]),.b(hsu[46]),.cin(hca[45]),.sum(fsu[674]),.carry(fca[674]));
FA FA675 (.a(fsu[531]),.b(fca[529]),.cin(fsu[532]),.sum(fsu[675]),.carry(fca[675]));
FA FA676 (.a(fca[530]),.b(fsu[533]),.cin(hca[46]),.sum(fsu[676]),.carry(fca[676]));
FA FA677 (.a(fsu[534]),.b(fca[531]),.cin(fsu[535]),.sum(fsu[677]),.carry(fca[677]));
FA FA678 (.a(fca[532]),.b(fsu[536]),.cin(fca[533]),.sum(fsu[678]),.carry(fca[678]));
FA FA679 (.a(fsu[537]),.b(fca[534]),.cin(fsu[538]),.sum(fsu[679]),.carry(fca[679]));
FA FA680 (.a(fca[535]),.b(fsu[539]),.cin(fca[536]),.sum(fsu[680]),.carry(fca[680]));
FA FA681 (.a(fsu[540]),.b(fca[537]),.cin(fsu[541]),.sum(fsu[681]),.carry(fca[681]));
FA FA682 (.a(fca[538]),.b(fsu[542]),.cin(fca[539]),.sum(fsu[682]),.carry(fca[682]));
FA FA683 (.a(fsu[543]),.b(fca[540]),.cin(fsu[544]),.sum(fsu[683]),.carry(fca[683]));
FA FA684 (.a(fca[541]),.b(fsu[545]),.cin(fca[542]),.sum(fsu[684]),.carry(fca[684]));
FA FA685 (.a(fsu[546]),.b(fca[543]),.cin(fsu[547]),.sum(fsu[685]),.carry(fca[685]));
FA FA686 (.a(fca[544]),.b(fsu[548]),.cin(fca[545]),.sum(fsu[686]),.carry(fca[686]));
FA FA687 (.a(fsu[549]),.b(fca[546]),.cin(fsu[550]),.sum(fsu[687]),.carry(fca[687]));
FA FA688 (.a(fca[547]),.b(fsu[551]),.cin(fca[548]),.sum(fsu[688]),.carry(fca[688]));
HA HA65 (.a(hsu[48]),.b(hca[47]),.sum_h(hsu[65]),.carry_h(hca[65]));
FA FA689 (.a(fsu[552]),.b(fca[549]),.cin(fsu[553]),.sum(fsu[689]),.carry(fca[689]));
FA FA690 (.a(fca[550]),.b(fsu[554]),.cin(fca[551]),.sum(fsu[690]),.carry(fca[690]));
HA HA66 (.a(fsu[555]),.b(hca[48]),.sum_h(hsu[66]),.carry_h(hca[66]));
FA FA691 (.a(fsu[556]),.b(fca[552]),.cin(fsu[557]),.sum(fsu[691]),.carry(fca[691]));
FA FA692 (.a(fca[553]),.b(fsu[558]),.cin(fca[554]),.sum(fsu[692]),.carry(fca[692]));
HA HA67 (.a(fsu[559]),.b(fca[555]),.sum_h(hsu[67]),.carry_h(hca[67]));
FA FA693 (.a(fsu[560]),.b(fca[556]),.cin(fsu[561]),.sum(fsu[693]),.carry(fca[693]));
FA FA694 (.a(fca[557]),.b(fsu[562]),.cin(fca[558]),.sum(fsu[694]),.carry(fca[694]));
FA FA695 (.a(fsu[563]),.b(fca[559]),.cin(pp[0][27]),.sum(fsu[695]),.carry(fca[695]));
FA FA696 (.a(fsu[564]),.b(fca[560]),.cin(fsu[565]),.sum(fsu[696]),.carry(fca[696]));
FA FA697 (.a(fca[561]),.b(fsu[566]),.cin(fca[562]),.sum(fsu[697]),.carry(fca[697]));
FA FA698 (.a(fsu[567]),.b(fca[563]),.cin(hsu[10]),.sum(fsu[698]),.carry(fca[698]));
FA FA699 (.a(fsu[568]),.b(fca[564]),.cin(fsu[569]),.sum(fsu[699]),.carry(fca[699]));
FA FA700 (.a(fca[565]),.b(fsu[570]),.cin(fca[566]),.sum(fsu[700]),.carry(fca[700]));
FA FA701 (.a(fsu[571]),.b(fca[567]),.cin(hsu[30]),.sum(fsu[701]),.carry(fca[701]));
FA FA702 (.a(fsu[572]),.b(fca[568]),.cin(fsu[573]),.sum(fsu[702]),.carry(fca[702]));
FA FA703 (.a(fca[569]),.b(fsu[574]),.cin(fca[570]),.sum(fsu[703]),.carry(fca[703]));
FA FA704 (.a(fsu[575]),.b(fca[571]),.cin(hsu[49]),.sum(fsu[704]),.carry(fca[704]));
FA FA705 (.a(fsu[576]),.b(fca[572]),.cin(fsu[577]),.sum(fsu[705]),.carry(fca[705]));
FA FA706 (.a(fca[573]),.b(fsu[578]),.cin(fca[574]),.sum(fsu[706]),.carry(fca[706]));
FA FA707 (.a(fsu[579]),.b(fca[575]),.cin(fsu[580]),.sum(fsu[707]),.carry(fca[707]));
FA FA708 (.a(fsu[581]),.b(fca[576]),.cin(fsu[582]),.sum(fsu[708]),.carry(fca[708]));
FA FA709 (.a(fca[577]),.b(fsu[583]),.cin(fca[578]),.sum(fsu[709]),.carry(fca[709]));
FA FA710 (.a(fsu[584]),.b(fca[579]),.cin(fsu[585]),.sum(fsu[710]),.carry(fca[710]));
FA FA711 (.a(fsu[586]),.b(fca[581]),.cin(fsu[587]),.sum(fsu[711]),.carry(fca[711]));
FA FA712 (.a(fca[582]),.b(fsu[588]),.cin(fca[583]),.sum(fsu[712]),.carry(fca[712]));
FA FA713 (.a(fsu[589]),.b(fca[584]),.cin(fsu[590]),.sum(fsu[713]),.carry(fca[713]));
FA FA714 (.a(fsu[591]),.b(fca[586]),.cin(fsu[592]),.sum(fsu[714]),.carry(fca[714]));
FA FA715 (.a(fca[587]),.b(fsu[593]),.cin(fca[588]),.sum(fsu[715]),.carry(fca[715]));
FA FA716 (.a(fsu[594]),.b(fca[589]),.cin(fsu[595]),.sum(fsu[716]),.carry(fca[716]));
FA FA717 (.a(hsu[50]),.b(fca[591]),.cin(fsu[596]),.sum(fsu[717]),.carry(fca[717]));
FA FA718 (.a(fca[592]),.b(fsu[597]),.cin(fca[593]),.sum(fsu[718]),.carry(fca[718]));
FA FA719 (.a(fsu[598]),.b(fca[594]),.cin(fsu[599]),.sum(fsu[719]),.carry(fca[719]));
FA FA720 (.a(hsu[51]),.b(hca[50]),.cin(fsu[600]),.sum(fsu[720]),.carry(fca[720]));
FA FA721 (.a(fca[596]),.b(fsu[601]),.cin(fca[597]),.sum(fsu[721]),.carry(fca[721]));
FA FA722 (.a(fsu[602]),.b(fca[598]),.cin(fsu[603]),.sum(fsu[722]),.carry(fca[722]));
FA FA723 (.a(hsu[31]),.b(hca[51]),.cin(fsu[604]),.sum(fsu[723]),.carry(fca[723]));
FA FA724 (.a(fca[600]),.b(fsu[605]),.cin(fca[601]),.sum(fsu[724]),.carry(fca[724]));
FA FA725 (.a(fsu[606]),.b(fca[602]),.cin(fsu[607]),.sum(fsu[725]),.carry(fca[725]));
HA HA68 (.a(hsu[32]),.b(fsu[608]),.sum_h(hsu[68]),.carry_h(hca[68]));
FA FA726 (.a(fca[604]),.b(fsu[609]),.cin(fca[605]),.sum(fsu[726]),.carry(fca[726]));
FA FA727 (.a(fsu[610]),.b(fca[606]),.cin(fsu[611]),.sum(fsu[727]),.carry(fca[727]));
HA HA69 (.a(hsu[33]),.b(fsu[612]),.sum_h(hsu[69]),.carry_h(hca[69]));
FA FA728 (.a(fca[608]),.b(fsu[613]),.cin(fca[609]),.sum(fsu[728]),.carry(fca[728]));
FA FA729 (.a(fsu[614]),.b(fca[610]),.cin(fsu[615]),.sum(fsu[729]),.carry(fca[729]));
FA FA730 (.a(fca[612]),.b(fsu[617]),.cin(fca[613]),.sum(fsu[730]),.carry(fca[730]));
FA FA731 (.a(fsu[618]),.b(fca[614]),.cin(fsu[619]),.sum(fsu[731]),.carry(fca[731]));
FA FA732 (.a(fca[616]),.b(fsu[620]),.cin(fca[617]),.sum(fsu[732]),.carry(fca[732]));
FA FA733 (.a(fsu[621]),.b(fca[618]),.cin(fsu[622]),.sum(fsu[733]),.carry(fca[733]));
FA FA734 (.a(hca[52]),.b(fsu[623]),.cin(fca[620]),.sum(fsu[734]),.carry(fca[734]));
FA FA735 (.a(fsu[624]),.b(fca[621]),.cin(fsu[625]),.sum(fsu[735]),.carry(fca[735]));
FA FA736 (.a(hca[53]),.b(fsu[626]),.cin(fca[623]),.sum(fsu[736]),.carry(fca[736]));
FA FA737 (.a(fsu[627]),.b(fca[624]),.cin(fsu[628]),.sum(fsu[737]),.carry(fca[737]));
FA FA738 (.a(hca[54]),.b(fsu[629]),.cin(fca[626]),.sum(fsu[738]),.carry(fca[738]));
FA FA739 (.a(fsu[630]),.b(fca[627]),.cin(fsu[631]),.sum(fsu[739]),.carry(fca[739]));
FA FA740 (.a(pp[31][14]),.b(fsu[632]),.cin(fca[629]),.sum(fsu[740]),.carry(fca[740]));
FA FA741 (.a(fsu[633]),.b(fca[630]),.cin(fsu[634]),.sum(fsu[741]),.carry(fca[741]));
HA HA70 (.a(fsu[635]),.b(fca[632]),.sum_h(hsu[70]),.carry_h(hca[70]));
FA FA742 (.a(fsu[636]),.b(fca[633]),.cin(fsu[637]),.sum(fsu[742]),.carry(fca[742]));
HA HA71 (.a(fsu[638]),.b(fca[635]),.sum_h(hsu[71]),.carry_h(hca[71]));
FA FA743 (.a(fsu[639]),.b(fca[636]),.cin(fsu[640]),.sum(fsu[743]),.carry(fca[743]));
HA HA72 (.a(fsu[641]),.b(fca[638]),.sum_h(hsu[72]),.carry_h(hca[72]));
FA FA744 (.a(fsu[642]),.b(fca[639]),.cin(fsu[643]),.sum(fsu[744]),.carry(fca[744]));
HA HA73 (.a(hsu[55]),.b(fca[641]),.sum_h(hsu[73]),.carry_h(hca[73]));
FA FA745 (.a(fsu[644]),.b(fca[642]),.cin(fsu[645]),.sum(fsu[745]),.carry(fca[745]));
HA HA74 (.a(fsu[494]),.b(hca[55]),.sum_h(hsu[74]),.carry_h(hca[74]));
FA FA746 (.a(fsu[646]),.b(fca[644]),.cin(fsu[647]),.sum(fsu[746]),.carry(fca[746]));
FA FA747 (.a(fsu[648]),.b(fca[646]),.cin(fsu[649]),.sum(fsu[747]),.carry(fca[747]));
FA FA748 (.a(fsu[650]),.b(fca[648]),.cin(fsu[651]),.sum(fsu[748]),.carry(fca[748]));
FA FA749 (.a(fsu[652]),.b(fca[650]),.cin(fsu[653]),.sum(fsu[749]),.carry(fca[749]));
FA FA750 (.a(fsu[654]),.b(fca[652]),.cin(fsu[655]),.sum(fsu[750]),.carry(fca[750]));
FA FA751 (.a(hsu[56]),.b(fca[654]),.cin(fsu[656]),.sum(fsu[751]),.carry(fca[751]));
FA FA752 (.a(hsu[57]),.b(hca[56]),.cin(fsu[657]),.sum(fsu[752]),.carry(fca[752]));
FA FA753 (.a(hsu[58]),.b(hca[57]),.cin(fsu[658]),.sum(fsu[753]),.carry(fca[753]));
FA FA754 (.a(hca[39]),.b(hca[58]),.cin(fsu[659]),.sum(fsu[754]),.carry(fca[754]));
//5th stage
HA HA75 (.a(hsu[60]),.b(hca[59]),.sum_h(z[5]),.carry_h(hca[75]));
HA HA76 (.a(hsu[61]),.b(hca[60]),.sum_h(hsu[76]),.carry_h(hca[76]));
HA HA77 (.a(fsu[663]),.b(hca[61]),.sum_h(hsu[77]),.carry_h(hca[77]));
HA HA78 (.a(fsu[664]),.b(fca[663]),.sum_h(hsu[78]),.carry_h(hca[78]));
HA HA79 (.a(fsu[665]),.b(fca[664]),.sum_h(hsu[79]),.carry_h(hca[79]));
FA FA755 (.a(fsu[666]),.b(fca[665]),.cin(hca[42]),.sum(fsu[755]),.carry(fca[755]));
FA FA756 (.a(fsu[667]),.b(fca[666]),.cin(hca[43]),.sum(fsu[756]),.carry(fca[756]));
FA FA757 (.a(fsu[668]),.b(fca[667]),.cin(hca[44]),.sum(fsu[757]),.carry(fca[757]));
FA FA758 (.a(fsu[669]),.b(fca[668]),.cin(fca[520]),.sum(fsu[758]),.carry(fca[758]));
FA FA759 (.a(fsu[670]),.b(fca[669]),.cin(hsu[62]),.sum(fsu[759]),.carry(fca[759]));
FA FA760 (.a(fsu[671]),.b(fca[670]),.cin(hsu[63]),.sum(fsu[760]),.carry(fca[760]));
FA FA761 (.a(fsu[672]),.b(fca[671]),.cin(hsu[64]),.sum(fsu[761]),.carry(fca[761]));
FA FA762 (.a(fsu[673]),.b(fca[672]),.cin(fsu[674]),.sum(fsu[762]),.carry(fca[762]));
FA FA763 (.a(fsu[675]),.b(fca[673]),.cin(fsu[676]),.sum(fsu[763]),.carry(fca[763]));
FA FA764 (.a(fsu[677]),.b(fca[675]),.cin(fsu[678]),.sum(fsu[764]),.carry(fca[764]));
FA FA765 (.a(fsu[679]),.b(fca[677]),.cin(fsu[680]),.sum(fsu[765]),.carry(fca[765]));
FA FA766 (.a(fsu[681]),.b(fca[679]),.cin(fsu[682]),.sum(fsu[766]),.carry(fca[766]));
HA HA80 (.a(fca[680]),.b(hca[27]),.sum_h(hsu[80]),.carry_h(hca[80]));
FA FA767 (.a(fsu[683]),.b(fca[681]),.cin(fsu[684]),.sum(fsu[767]),.carry(fca[767]));
HA HA81 (.a(fca[682]),.b(fca[349]),.sum_h(hsu[81]),.carry_h(hca[81]));
FA FA768 (.a(fsu[685]),.b(fca[683]),.cin(fsu[686]),.sum(fsu[768]),.carry(fca[768]));
HA HA82 (.a(fca[684]),.b(hsu[47]),.sum_h(hsu[82]),.carry_h(hca[82]));
FA FA769 (.a(fsu[687]),.b(fca[685]),.cin(fsu[688]),.sum(fsu[769]),.carry(fca[769]));
HA HA83 (.a(fca[686]),.b(hsu[65]),.sum_h(hsu[83]),.carry_h(hca[83]));
FA FA770 (.a(fsu[689]),.b(fca[687]),.cin(fsu[690]),.sum(fsu[770]),.carry(fca[770]));
FA FA771 (.a(fca[688]),.b(hsu[66]),.cin(hca[65]),.sum(fsu[771]),.carry(fca[771]));
FA FA772 (.a(fsu[691]),.b(fca[689]),.cin(fsu[692]),.sum(fsu[772]),.carry(fca[772]));
FA FA773 (.a(fca[690]),.b(hsu[67]),.cin(hca[66]),.sum(fsu[773]),.carry(fca[773]));
FA FA774 (.a(fsu[693]),.b(fca[691]),.cin(fsu[694]),.sum(fsu[774]),.carry(fca[774]));
FA FA775 (.a(fca[692]),.b(fsu[695]),.cin(hca[67]),.sum(fsu[775]),.carry(fca[775]));
FA FA776 (.a(fsu[696]),.b(fca[693]),.cin(fsu[697]),.sum(fsu[776]),.carry(fca[776]));
FA FA777 (.a(fca[694]),.b(fsu[698]),.cin(fca[695]),.sum(fsu[777]),.carry(fca[777]));
FA FA778 (.a(fsu[699]),.b(fca[696]),.cin(fsu[700]),.sum(fsu[778]),.carry(fca[778]));
FA FA779 (.a(fca[697]),.b(fsu[701]),.cin(fca[698]),.sum(fsu[779]),.carry(fca[779]));
FA FA780 (.a(fsu[702]),.b(fca[699]),.cin(fsu[703]),.sum(fsu[780]),.carry(fca[780]));
FA FA781 (.a(fca[700]),.b(fsu[704]),.cin(fca[701]),.sum(fsu[781]),.carry(fca[781]));
FA FA782 (.a(fsu[705]),.b(fca[702]),.cin(fsu[706]),.sum(fsu[782]),.carry(fca[782]));
FA FA783 (.a(fca[703]),.b(fsu[707]),.cin(fca[704]),.sum(fsu[783]),.carry(fca[783]));
FA FA784 (.a(fsu[708]),.b(fca[705]),.cin(fsu[709]),.sum(fsu[784]),.carry(fca[784]));
FA FA785 (.a(fca[706]),.b(fsu[710]),.cin(fca[707]),.sum(fsu[785]),.carry(fca[785]));
FA FA786 (.a(fsu[711]),.b(fca[708]),.cin(fsu[712]),.sum(fsu[786]),.carry(fca[786]));
FA FA787 (.a(fca[709]),.b(fsu[713]),.cin(fca[710]),.sum(fsu[787]),.carry(fca[787]));
FA FA788 (.a(fsu[714]),.b(fca[711]),.cin(fsu[715]),.sum(fsu[788]),.carry(fca[788]));
FA FA789 (.a(fca[712]),.b(fsu[716]),.cin(fca[713]),.sum(fsu[789]),.carry(fca[789]));
FA FA790 (.a(fsu[717]),.b(fca[714]),.cin(fsu[718]),.sum(fsu[790]),.carry(fca[790]));
FA FA791 (.a(fca[715]),.b(fsu[719]),.cin(fca[716]),.sum(fsu[791]),.carry(fca[791]));
FA FA792 (.a(fsu[720]),.b(fca[717]),.cin(fsu[721]),.sum(fsu[792]),.carry(fca[792]));
FA FA793 (.a(fca[718]),.b(fsu[722]),.cin(fca[719]),.sum(fsu[793]),.carry(fca[793]));
FA FA794 (.a(fsu[723]),.b(fca[720]),.cin(fsu[724]),.sum(fsu[794]),.carry(fca[794]));
FA FA795 (.a(fca[721]),.b(fsu[725]),.cin(fca[722]),.sum(fsu[795]),.carry(fca[795]));
FA FA796 (.a(hsu[68]),.b(fca[723]),.cin(fsu[726]),.sum(fsu[796]),.carry(fca[796]));
FA FA797 (.a(fca[724]),.b(fsu[727]),.cin(fca[725]),.sum(fsu[797]),.carry(fca[797]));
FA FA798 (.a(hsu[69]),.b(hca[68]),.cin(fsu[728]),.sum(fsu[798]),.carry(fca[798]));
FA FA799 (.a(fca[726]),.b(fsu[729]),.cin(fca[727]),.sum(fsu[799]),.carry(fca[799]));
FA FA800 (.a(fsu[616]),.b(hca[69]),.cin(fsu[730]),.sum(fsu[800]),.carry(fca[800]));
FA FA801 (.a(fca[728]),.b(fsu[731]),.cin(fca[729]),.sum(fsu[801]),.carry(fca[801]));
HA HA84 (.a(hsu[52]),.b(fsu[732]),.sum_h(hsu[84]),.carry_h(hca[84]));
FA FA802 (.a(fca[730]),.b(fsu[733]),.cin(fca[731]),.sum(fsu[802]),.carry(fca[802]));
HA HA85 (.a(hsu[53]),.b(fsu[734]),.sum_h(hsu[85]),.carry_h(hca[85]));
FA FA803 (.a(fca[732]),.b(fsu[735]),.cin(fca[733]),.sum(fsu[803]),.carry(fca[803]));
HA HA86 (.a(hsu[54]),.b(fsu[736]),.sum_h(hsu[86]),.carry_h(hca[86]));
FA FA804 (.a(fca[734]),.b(fsu[737]),.cin(fca[735]),.sum(fsu[804]),.carry(fca[804]));
HA HA87 (.a(hsu[15]),.b(fsu[738]),.sum_h(hsu[87]),.carry_h(hca[87]));
FA FA805 (.a(fca[736]),.b(fsu[739]),.cin(fca[737]),.sum(fsu[805]),.carry(fca[805]));
FA FA806 (.a(fca[738]),.b(fsu[741]),.cin(fca[739]),.sum(fsu[806]),.carry(fca[806]));
FA FA807 (.a(fca[740]),.b(fsu[742]),.cin(fca[741]),.sum(fsu[807]),.carry(fca[807]));
FA FA808 (.a(hca[70]),.b(fsu[743]),.cin(fca[742]),.sum(fsu[808]),.carry(fca[808]));
FA FA809 (.a(hca[71]),.b(fsu[744]),.cin(fca[743]),.sum(fsu[809]),.carry(fca[809]));
FA FA810 (.a(hca[72]),.b(fsu[745]),.cin(fca[744]),.sum(fsu[810]),.carry(fca[810]));
FA FA811 (.a(hca[73]),.b(fsu[746]),.cin(fca[745]),.sum(fsu[811]),.carry(fca[811]));
FA FA812 (.a(hca[74]),.b(fsu[747]),.cin(fca[746]),.sum(fsu[812]),.carry(fca[812]));
FA FA813 (.a(fsu[289]),.b(fsu[748]),.cin(fca[747]),.sum(fsu[813]),.carry(fca[813]));
HA HA88 (.a(fsu[749]),.b(fca[748]),.sum_h(hsu[88]),.carry_h(hca[88]));
HA HA89 (.a(fsu[750]),.b(fca[749]),.sum_h(hsu[89]),.carry_h(hca[89]));
HA HA90 (.a(fsu[751]),.b(fca[750]),.sum_h(hsu[90]),.carry_h(hca[90]));
HA HA91 (.a(fsu[752]),.b(fca[751]),.sum_h(hsu[91]),.carry_h(hca[91]));
HA HA92 (.a(fsu[753]),.b(fca[752]),.sum_h(hsu[92]),.carry_h(hca[92]));
HA HA93 (.a(fsu[754]),.b(fca[753]),.sum_h(hsu[93]),.carry_h(hca[93]));
HA HA94 (.a(fsu[660]),.b(fca[754]),.sum_h(hsu[94]),.carry_h(hca[94]));
//6th stage
HA HA95 (.a(hsu[76]),.b(hca[75]),.sum_h(z[6]),.carry_h(hca[95]));
HA HA96 (.a(hsu[77]),.b(hca[76]),.sum_h(hsu[96]),.carry_h(hca[96]));
HA HA97 (.a(hsu[78]),.b(hca[77]),.sum_h(hsu[97]),.carry_h(hca[97]));
HA HA98 (.a(hsu[79]),.b(hca[78]),.sum_h(hsu[98]),.carry_h(hca[98]));
HA HA99 (.a(fsu[755]),.b(hca[79]),.sum_h(hsu[99]),.carry_h(hca[99]));
HA HA100 (.a(fsu[756]),.b(fca[755]),.sum_h(hsu[100]),.carry_h(hca[100]));
HA HA101 (.a(fsu[757]),.b(fca[756]),.sum_h(hsu[101]),.carry_h(hca[101]));
HA HA102 (.a(fsu[758]),.b(fca[757]),.sum_h(hsu[102]),.carry_h(hca[102]));
HA HA103 (.a(fsu[759]),.b(fca[758]),.sum_h(hsu[103]),.carry_h(hca[103]));
FA FA814 (.a(fsu[760]),.b(fca[759]),.cin(hca[62]),.sum(fsu[814]),.carry(fca[814]));
FA FA815 (.a(fsu[761]),.b(fca[760]),.cin(hca[63]),.sum(fsu[815]),.carry(fca[815]));
FA FA816 (.a(fsu[762]),.b(fca[761]),.cin(hca[64]),.sum(fsu[816]),.carry(fca[816]));
FA FA817 (.a(fsu[763]),.b(fca[762]),.cin(fca[674]),.sum(fsu[817]),.carry(fca[817]));
FA FA818 (.a(fsu[764]),.b(fca[763]),.cin(fca[676]),.sum(fsu[818]),.carry(fca[818]));
FA FA819 (.a(fsu[765]),.b(fca[764]),.cin(fca[678]),.sum(fsu[819]),.carry(fca[819]));
FA FA820 (.a(fsu[766]),.b(fca[765]),.cin(hsu[80]),.sum(fsu[820]),.carry(fca[820]));
FA FA821 (.a(fsu[767]),.b(fca[766]),.cin(hsu[81]),.sum(fsu[821]),.carry(fca[821]));
FA FA822 (.a(fsu[768]),.b(fca[767]),.cin(hsu[82]),.sum(fsu[822]),.carry(fca[822]));
FA FA823 (.a(fsu[769]),.b(fca[768]),.cin(hsu[83]),.sum(fsu[823]),.carry(fca[823]));
FA FA824 (.a(fsu[770]),.b(fca[769]),.cin(fsu[771]),.sum(fsu[824]),.carry(fca[824]));
FA FA825 (.a(fsu[772]),.b(fca[770]),.cin(fsu[773]),.sum(fsu[825]),.carry(fca[825]));
FA FA826 (.a(fsu[774]),.b(fca[772]),.cin(fsu[775]),.sum(fsu[826]),.carry(fca[826]));
FA FA827 (.a(fsu[776]),.b(fca[774]),.cin(fsu[777]),.sum(fsu[827]),.carry(fca[827]));
FA FA828 (.a(fsu[778]),.b(fca[776]),.cin(fsu[779]),.sum(fsu[828]),.carry(fca[828]));
FA FA829 (.a(fsu[780]),.b(fca[778]),.cin(fsu[781]),.sum(fsu[829]),.carry(fca[829]));
FA FA830 (.a(fsu[782]),.b(fca[780]),.cin(fsu[783]),.sum(fsu[830]),.carry(fca[830]));
FA FA831 (.a(fsu[784]),.b(fca[782]),.cin(fsu[785]),.sum(fsu[831]),.carry(fca[831]));
FA FA832 (.a(fsu[786]),.b(fca[784]),.cin(fsu[787]),.sum(fsu[832]),.carry(fca[832]));
FA FA833 (.a(fsu[788]),.b(fca[786]),.cin(fsu[789]),.sum(fsu[833]),.carry(fca[833]));
FA FA834 (.a(fsu[790]),.b(fca[788]),.cin(fsu[791]),.sum(fsu[834]),.carry(fca[834]));
FA FA835 (.a(fsu[792]),.b(fca[790]),.cin(fsu[793]),.sum(fsu[835]),.carry(fca[835]));
FA FA836 (.a(fsu[794]),.b(fca[792]),.cin(fsu[795]),.sum(fsu[836]),.carry(fca[836]));
FA FA837 (.a(fsu[796]),.b(fca[794]),.cin(fsu[797]),.sum(fsu[837]),.carry(fca[837]));
FA FA838 (.a(fsu[798]),.b(fca[796]),.cin(fsu[799]),.sum(fsu[838]),.carry(fca[838]));
FA FA839 (.a(fsu[800]),.b(fca[798]),.cin(fsu[801]),.sum(fsu[839]),.carry(fca[839]));
FA FA840 (.a(hsu[84]),.b(fca[800]),.cin(fsu[802]),.sum(fsu[840]),.carry(fca[840]));
FA FA841 (.a(hsu[85]),.b(hca[84]),.cin(fsu[803]),.sum(fsu[841]),.carry(fca[841]));
FA FA842 (.a(hsu[86]),.b(hca[85]),.cin(fsu[804]),.sum(fsu[842]),.carry(fca[842]));
FA FA843 (.a(hsu[87]),.b(hca[86]),.cin(fsu[805]),.sum(fsu[843]),.carry(fca[843]));
FA FA844 (.a(fsu[740]),.b(hca[87]),.cin(fsu[806]),.sum(fsu[844]),.carry(fca[844]));
HA HA104 (.a(hsu[70]),.b(fsu[807]),.sum_h(hsu[104]),.carry_h(hca[104]));
HA HA105 (.a(hsu[71]),.b(fsu[808]),.sum_h(hsu[105]),.carry_h(hca[105]));
HA HA106 (.a(hsu[72]),.b(fsu[809]),.sum_h(hsu[106]),.carry_h(hca[106]));
HA HA107 (.a(hsu[73]),.b(fsu[810]),.sum_h(hsu[107]),.carry_h(hca[107]));
HA HA108 (.a(hsu[74]),.b(fsu[811]),.sum_h(hsu[108]),.carry_h(hca[108]));
HA HA109 (.a(fsu[497]),.b(fsu[812]),.sum_h(hsu[109]),.carry_h(hca[109]));
//7th stage
HA HA110 (.a(hsu[96]),.b(hca[95]),.sum_h(z[7]),.carry_h(hca[110]));
HA HA111 (.a(hsu[97]),.b(hca[96]),.sum_h(hsu[111]),.carry_h(hca[111]));
HA HA112 (.a(hsu[98]),.b(hca[97]),.sum_h(hsu[112]),.carry_h(hca[112]));
HA HA113 (.a(hsu[99]),.b(hca[98]),.sum_h(hsu[113]),.carry_h(hca[113]));
HA HA114 (.a(hsu[100]),.b(hca[99]),.sum_h(hsu[114]),.carry_h(hca[114]));
HA HA115 (.a(hsu[101]),.b(hca[100]),.sum_h(hsu[115]),.carry_h(hca[115]));
HA HA116 (.a(hsu[102]),.b(hca[101]),.sum_h(hsu[116]),.carry_h(hca[116]));
HA HA117 (.a(hsu[103]),.b(hca[102]),.sum_h(hsu[117]),.carry_h(hca[117]));
HA HA118 (.a(fsu[814]),.b(hca[103]),.sum_h(hsu[118]),.carry_h(hca[118]));
HA HA119 (.a(fsu[815]),.b(fca[814]),.sum_h(hsu[119]),.carry_h(hca[119]));
HA HA120 (.a(fsu[816]),.b(fca[815]),.sum_h(hsu[120]),.carry_h(hca[120]));
HA HA121 (.a(fsu[817]),.b(fca[816]),.sum_h(hsu[121]),.carry_h(hca[121]));
HA HA122 (.a(fsu[818]),.b(fca[817]),.sum_h(hsu[122]),.carry_h(hca[122]));
HA HA123 (.a(fsu[819]),.b(fca[818]),.sum_h(hsu[123]),.carry_h(hca[123]));
HA HA124 (.a(fsu[820]),.b(fca[819]),.sum_h(hsu[124]),.carry_h(hca[124]));
FA FA845 (.a(fsu[821]),.b(fca[820]),.cin(hca[80]),.sum(fsu[845]),.carry(fca[845]));
FA FA846 (.a(fsu[822]),.b(fca[821]),.cin(hca[81]),.sum(fsu[846]),.carry(fca[846]));
FA FA847 (.a(fsu[823]),.b(fca[822]),.cin(hca[82]),.sum(fsu[847]),.carry(fca[847]));
FA FA848 (.a(fsu[824]),.b(fca[823]),.cin(hca[83]),.sum(fsu[848]),.carry(fca[848]));
FA FA849 (.a(fsu[825]),.b(fca[824]),.cin(fca[771]),.sum(fsu[849]),.carry(fca[849]));
FA FA850 (.a(fsu[826]),.b(fca[825]),.cin(fca[773]),.sum(fsu[850]),.carry(fca[850]));
FA FA851 (.a(fsu[827]),.b(fca[826]),.cin(fca[775]),.sum(fsu[851]),.carry(fca[851]));
FA FA852 (.a(fsu[828]),.b(fca[827]),.cin(fca[777]),.sum(fsu[852]),.carry(fca[852]));
FA FA853 (.a(fsu[829]),.b(fca[828]),.cin(fca[779]),.sum(fsu[853]),.carry(fca[853]));
FA FA854 (.a(fsu[830]),.b(fca[829]),.cin(fca[781]),.sum(fsu[854]),.carry(fca[854]));
FA FA855 (.a(fsu[831]),.b(fca[830]),.cin(fca[783]),.sum(fsu[855]),.carry(fca[855]));
FA FA856 (.a(fsu[832]),.b(fca[831]),.cin(fca[785]),.sum(fsu[856]),.carry(fca[856]));
FA FA857 (.a(fsu[833]),.b(fca[832]),.cin(fca[787]),.sum(fsu[857]),.carry(fca[857]));
FA FA858 (.a(fsu[834]),.b(fca[833]),.cin(fca[789]),.sum(fsu[858]),.carry(fca[858]));
FA FA859 (.a(fsu[835]),.b(fca[834]),.cin(fca[791]),.sum(fsu[859]),.carry(fca[859]));
FA FA860 (.a(fsu[836]),.b(fca[835]),.cin(fca[793]),.sum(fsu[860]),.carry(fca[860]));
FA FA861 (.a(fsu[837]),.b(fca[836]),.cin(fca[795]),.sum(fsu[861]),.carry(fca[861]));
FA FA862 (.a(fsu[838]),.b(fca[837]),.cin(fca[797]),.sum(fsu[862]),.carry(fca[862]));
FA FA863 (.a(fsu[839]),.b(fca[838]),.cin(fca[799]),.sum(fsu[863]),.carry(fca[863]));
FA FA864 (.a(fsu[840]),.b(fca[839]),.cin(fca[801]),.sum(fsu[864]),.carry(fca[864]));
FA FA865 (.a(fsu[841]),.b(fca[840]),.cin(fca[802]),.sum(fsu[865]),.carry(fca[865]));
FA FA866 (.a(fsu[842]),.b(fca[841]),.cin(fca[803]),.sum(fsu[866]),.carry(fca[866]));
FA FA867 (.a(fsu[843]),.b(fca[842]),.cin(fca[804]),.sum(fsu[867]),.carry(fca[867]));
FA FA868 (.a(fsu[844]),.b(fca[843]),.cin(fca[805]),.sum(fsu[868]),.carry(fca[868]));
FA FA869 (.a(hsu[104]),.b(fca[844]),.cin(fca[806]),.sum(fsu[869]),.carry(fca[869]));
FA FA870 (.a(hsu[105]),.b(hca[104]),.cin(fca[807]),.sum(fsu[870]),.carry(fca[870]));
FA FA871 (.a(hsu[106]),.b(hca[105]),.cin(fca[808]),.sum(fsu[871]),.carry(fca[871]));
FA FA872 (.a(hsu[107]),.b(hca[106]),.cin(fca[809]),.sum(fsu[872]),.carry(fca[872]));
FA FA873 (.a(hsu[108]),.b(hca[107]),.cin(fca[810]),.sum(fsu[873]),.carry(fca[873]));
FA FA874 (.a(hsu[109]),.b(hca[108]),.cin(fca[811]),.sum(fsu[874]),.carry(fca[874]));
FA FA875 (.a(fsu[813]),.b(hca[109]),.cin(fca[812]),.sum(fsu[875]),.carry(fca[875]));
HA HA125 (.a(hsu[88]),.b(fca[813]),.sum_h(hsu[125]),.carry_h(hca[125]));
HA HA126 (.a(hsu[89]),.b(hca[88]),.sum_h(hsu[126]),.carry_h(hca[126]));
HA HA127 (.a(hsu[90]),.b(hca[89]),.sum_h(hsu[127]),.carry_h(hca[127]));
HA HA128 (.a(hsu[91]),.b(hca[90]),.sum_h(hsu[128]),.carry_h(hca[128]));
HA HA129 (.a(hsu[92]),.b(hca[91]),.sum_h(hsu[129]),.carry_h(hca[129]));
HA HA130 (.a(hsu[93]),.b(hca[92]),.sum_h(hsu[130]),.carry_h(hca[130]));
HA HA131 (.a(hsu[94]),.b(hca[93]),.sum_h(hsu[131]),.carry_h(hca[131]));
HA HA132 (.a(fsu[661]),.b(hca[94]),.sum_h(hsu[132]),.carry_h(hca[132]));
//8th stage
HA HA133 (.a(hsu[111]),.b(hca[110]),.sum_h(z[8]),.carry_h(hca[133]));
HA HA134 (.a(hsu[112]),.b(hca[111]),.sum_h(hsu[134]),.carry_h(hca[134]));
HA HA135 (.a(hsu[113]),.b(hca[112]),.sum_h(hsu[135]),.carry_h(hca[135]));
HA HA136 (.a(hsu[114]),.b(hca[113]),.sum_h(hsu[136]),.carry_h(hca[136]));
HA HA137 (.a(hsu[115]),.b(hca[114]),.sum_h(hsu[137]),.carry_h(hca[137]));
HA HA138 (.a(hsu[116]),.b(hca[115]),.sum_h(hsu[138]),.carry_h(hca[138]));
HA HA139 (.a(hsu[117]),.b(hca[116]),.sum_h(hsu[139]),.carry_h(hca[139]));
HA HA140 (.a(hsu[118]),.b(hca[117]),.sum_h(hsu[140]),.carry_h(hca[140]));
HA HA141 (.a(hsu[119]),.b(hca[118]),.sum_h(hsu[141]),.carry_h(hca[141]));
HA HA142 (.a(hsu[120]),.b(hca[119]),.sum_h(hsu[142]),.carry_h(hca[142]));
HA HA143 (.a(hsu[121]),.b(hca[120]),.sum_h(hsu[143]),.carry_h(hca[143]));
HA HA144 (.a(hsu[122]),.b(hca[121]),.sum_h(hsu[144]),.carry_h(hca[144]));
HA HA145 (.a(hsu[123]),.b(hca[122]),.sum_h(hsu[145]),.carry_h(hca[145]));
HA HA146 (.a(hsu[124]),.b(hca[123]),.sum_h(hsu[146]),.carry_h(hca[146]));
HA HA147 (.a(fsu[845]),.b(hca[124]),.sum_h(hsu[147]),.carry_h(hca[147]));
HA HA148 (.a(fsu[846]),.b(fca[845]),.sum_h(hsu[148]),.carry_h(hca[148]));
HA HA149 (.a(fsu[847]),.b(fca[846]),.sum_h(hsu[149]),.carry_h(hca[149]));
HA HA150 (.a(fsu[848]),.b(fca[847]),.sum_h(hsu[150]),.carry_h(hca[150]));
HA HA151 (.a(fsu[849]),.b(fca[848]),.sum_h(hsu[151]),.carry_h(hca[151]));
HA HA152 (.a(fsu[850]),.b(fca[849]),.sum_h(hsu[152]),.carry_h(hca[152]));
HA HA153 (.a(fsu[851]),.b(fca[850]),.sum_h(hsu[153]),.carry_h(hca[153]));
HA HA154 (.a(fsu[852]),.b(fca[851]),.sum_h(hsu[154]),.carry_h(hca[154]));
HA HA155 (.a(fsu[853]),.b(fca[852]),.sum_h(hsu[155]),.carry_h(hca[155]));
FA FA876 (.a(fsu[854]),.b(fca[853]),.cin(hca[49]),.sum(fsu[876]),.carry(fca[876]));
FA FA877 (.a(fsu[855]),.b(fca[854]),.cin(fca[580]),.sum(fsu[877]),.carry(fca[877]));
FA FA878 (.a(fsu[856]),.b(fca[855]),.cin(fca[585]),.sum(fsu[878]),.carry(fca[878]));
FA FA879 (.a(fsu[857]),.b(fca[856]),.cin(fca[590]),.sum(fsu[879]),.carry(fca[879]));
FA FA880 (.a(fsu[858]),.b(fca[857]),.cin(fca[595]),.sum(fsu[880]),.carry(fca[880]));
FA FA881 (.a(fsu[859]),.b(fca[858]),.cin(fca[599]),.sum(fsu[881]),.carry(fca[881]));
FA FA882 (.a(fsu[860]),.b(fca[859]),.cin(fca[603]),.sum(fsu[882]),.carry(fca[882]));
FA FA883 (.a(fsu[861]),.b(fca[860]),.cin(fca[607]),.sum(fsu[883]),.carry(fca[883]));
FA FA884 (.a(fsu[862]),.b(fca[861]),.cin(fca[611]),.sum(fsu[884]),.carry(fca[884]));
FA FA885 (.a(fsu[863]),.b(fca[862]),.cin(fca[615]),.sum(fsu[885]),.carry(fca[885]));
FA FA886 (.a(fsu[864]),.b(fca[863]),.cin(fca[619]),.sum(fsu[886]),.carry(fca[886]));
FA FA887 (.a(fsu[865]),.b(fca[864]),.cin(fca[622]),.sum(fsu[887]),.carry(fca[887]));
FA FA888 (.a(fsu[866]),.b(fca[865]),.cin(fca[625]),.sum(fsu[888]),.carry(fca[888]));
FA FA889 (.a(fsu[867]),.b(fca[866]),.cin(fca[628]),.sum(fsu[889]),.carry(fca[889]));
FA FA890 (.a(fsu[868]),.b(fca[867]),.cin(fca[631]),.sum(fsu[890]),.carry(fca[890]));
FA FA891 (.a(fsu[869]),.b(fca[868]),.cin(fca[634]),.sum(fsu[891]),.carry(fca[891]));
FA FA892 (.a(fsu[870]),.b(fca[869]),.cin(fca[637]),.sum(fsu[892]),.carry(fca[892]));
FA FA893 (.a(fsu[871]),.b(fca[870]),.cin(fca[640]),.sum(fsu[893]),.carry(fca[893]));
FA FA894 (.a(fsu[872]),.b(fca[871]),.cin(fca[643]),.sum(fsu[894]),.carry(fca[894]));
FA FA895 (.a(fsu[873]),.b(fca[872]),.cin(fca[645]),.sum(fsu[895]),.carry(fca[895]));
FA FA896 (.a(fsu[874]),.b(fca[873]),.cin(fca[647]),.sum(fsu[896]),.carry(fca[896]));
FA FA897 (.a(fsu[875]),.b(fca[874]),.cin(fca[649]),.sum(fsu[897]),.carry(fca[897]));
FA FA898 (.a(hsu[125]),.b(fca[875]),.cin(fca[651]),.sum(fsu[898]),.carry(fca[898]));
FA FA899 (.a(hsu[126]),.b(hca[125]),.cin(fca[653]),.sum(fsu[899]),.carry(fca[899]));
FA FA900 (.a(hsu[127]),.b(hca[126]),.cin(fca[655]),.sum(fsu[900]),.carry(fca[900]));
FA FA901 (.a(hsu[128]),.b(hca[127]),.cin(fca[656]),.sum(fsu[901]),.carry(fca[901]));
FA FA902 (.a(hsu[129]),.b(hca[128]),.cin(fca[657]),.sum(fsu[902]),.carry(fca[902]));
FA FA903 (.a(hsu[130]),.b(hca[129]),.cin(fca[658]),.sum(fsu[903]),.carry(fca[903]));
FA FA904 (.a(hsu[131]),.b(hca[130]),.cin(fca[659]),.sum(fsu[904]),.carry(fca[904]));
FA FA905 (.a(hsu[132]),.b(hca[131]),.cin(fca[660]),.sum(fsu[905]),.carry(fca[905]));
FA FA906 (.a(fsu[662]),.b(hca[132]),.cin(fca[661]),.sum(fsu[906]),.carry(fca[906]));
HA HA156 (.a(pp[31][31]),.b(fca[662]),.sum_h(hsu[156]),.carry_h(hca[156]));
//final
HA HA157 (.a(hsu[134]),.b(hca[133]),.sum_h(z[9]),.carry_h(hca[157]));
FA FA907 (.a(hsu[135]),.b(hca[134]),.cin(hca[157]),.sum(z[10]),.carry(fca[907]));
FA FA908 (.a(hsu[136]),.b(hca[135]),.cin(fca[907]),.sum(z[11]),.carry(fca[908]));
FA FA909 (.a(hsu[137]),.b(hca[136]),.cin(fca[908]),.sum(z[12]),.carry(fca[909]));
FA FA910 (.a(hsu[138]),.b(hca[137]),.cin(fca[909]),.sum(z[13]),.carry(fca[910]));
FA FA911 (.a(hsu[139]),.b(hca[138]),.cin(fca[910]),.sum(z[14]),.carry(fca[911]));
FA FA912 (.a(hsu[140]),.b(hca[139]),.cin(fca[911]),.sum(z[15]),.carry(fca[912]));
FA FA913 (.a(hsu[141]),.b(hca[140]),.cin(fca[912]),.sum(z[16]),.carry(fca[913]));
FA FA914 (.a(hsu[142]),.b(hca[141]),.cin(fca[913]),.sum(z[17]),.carry(fca[914]));
FA FA915 (.a(hsu[143]),.b(hca[142]),.cin(fca[914]),.sum(z[18]),.carry(fca[915]));
FA FA916 (.a(hsu[144]),.b(hca[143]),.cin(fca[915]),.sum(z[19]),.carry(fca[916]));
FA FA917 (.a(hsu[145]),.b(hca[144]),.cin(fca[916]),.sum(z[20]),.carry(fca[917]));
FA FA918 (.a(hsu[146]),.b(hca[145]),.cin(fca[917]),.sum(z[21]),.carry(fca[918]));
FA FA919 (.a(hsu[147]),.b(hca[146]),.cin(fca[918]),.sum(z[22]),.carry(fca[919]));
FA FA920 (.a(hsu[148]),.b(hca[147]),.cin(fca[919]),.sum(z[23]),.carry(fca[920]));
FA FA921 (.a(hsu[149]),.b(hca[148]),.cin(fca[920]),.sum(z[24]),.carry(fca[921]));
FA FA922 (.a(hsu[150]),.b(hca[149]),.cin(fca[921]),.sum(z[25]),.carry(fca[922]));
FA FA923 (.a(hsu[151]),.b(hca[150]),.cin(fca[922]),.sum(z[26]),.carry(fca[923]));
FA FA924 (.a(hsu[152]),.b(hca[151]),.cin(fca[923]),.sum(z[27]),.carry(fca[924]));
FA FA925 (.a(hsu[153]),.b(hca[152]),.cin(fca[924]),.sum(z[28]),.carry(fca[925]));
FA FA926 (.a(hsu[154]),.b(hca[153]),.cin(fca[925]),.sum(z[29]),.carry(fca[926]));
FA FA927 (.a(hsu[155]),.b(hca[154]),.cin(fca[926]),.sum(z[30]),.carry(fca[927]));
FA FA928 (.a(fsu[876]),.b(hca[155]),.cin(fca[927]),.sum(z[31]),.carry(fca[928]));
FA FA929 (.a(fsu[877]),.b(fca[876]),.cin(fca[928]),.sum(z[32]),.carry(fca[929]));
FA FA930 (.a(fsu[878]),.b(fca[877]),.cin(fca[929]),.sum(z[33]),.carry(fca[930]));
FA FA931 (.a(fsu[879]),.b(fca[878]),.cin(fca[930]),.sum(z[34]),.carry(fca[931]));
FA FA932 (.a(fsu[880]),.b(fca[879]),.cin(fca[931]),.sum(z[35]),.carry(fca[932]));
FA FA933 (.a(fsu[881]),.b(fca[880]),.cin(fca[932]),.sum(z[36]),.carry(fca[933]));
FA FA934 (.a(fsu[882]),.b(fca[881]),.cin(fca[933]),.sum(z[37]),.carry(fca[934]));
FA FA935 (.a(fsu[883]),.b(fca[882]),.cin(fca[934]),.sum(z[38]),.carry(fca[935]));
FA FA936 (.a(fsu[884]),.b(fca[883]),.cin(fca[935]),.sum(z[39]),.carry(fca[936]));
FA FA937 (.a(fsu[885]),.b(fca[884]),.cin(fca[936]),.sum(z[40]),.carry(fca[937]));
FA FA938 (.a(fsu[886]),.b(fca[885]),.cin(fca[937]),.sum(z[41]),.carry(fca[938]));
FA FA939 (.a(fsu[887]),.b(fca[886]),.cin(fca[938]),.sum(z[42]),.carry(fca[939]));
FA FA940 (.a(fsu[888]),.b(fca[887]),.cin(fca[939]),.sum(z[43]),.carry(fca[940]));
FA FA941 (.a(fsu[889]),.b(fca[888]),.cin(fca[940]),.sum(z[44]),.carry(fca[941]));
FA FA942 (.a(fsu[890]),.b(fca[889]),.cin(fca[941]),.sum(z[45]),.carry(fca[942]));
FA FA943 (.a(fsu[891]),.b(fca[890]),.cin(fca[942]),.sum(z[46]),.carry(fca[943]));
FA FA944 (.a(fsu[892]),.b(fca[891]),.cin(fca[943]),.sum(z[47]),.carry(fca[944]));
FA FA945 (.a(fsu[893]),.b(fca[892]),.cin(fca[944]),.sum(z[48]),.carry(fca[945]));
FA FA946 (.a(fsu[894]),.b(fca[893]),.cin(fca[945]),.sum(z[49]),.carry(fca[946]));
FA FA947 (.a(fsu[895]),.b(fca[894]),.cin(fca[946]),.sum(z[50]),.carry(fca[947]));
FA FA948 (.a(fsu[896]),.b(fca[895]),.cin(fca[947]),.sum(z[51]),.carry(fca[948]));
FA FA949 (.a(fsu[897]),.b(fca[896]),.cin(fca[948]),.sum(z[52]),.carry(fca[949]));
FA FA950 (.a(fsu[898]),.b(fca[897]),.cin(fca[949]),.sum(z[53]),.carry(fca[950]));
FA FA951 (.a(fsu[899]),.b(fca[898]),.cin(fca[950]),.sum(z[54]),.carry(fca[951]));
FA FA952 (.a(fsu[900]),.b(fca[899]),.cin(fca[951]),.sum(z[55]),.carry(fca[952]));
FA FA953 (.a(fsu[901]),.b(fca[900]),.cin(fca[952]),.sum(z[56]),.carry(fca[953]));
FA FA954 (.a(fsu[902]),.b(fca[901]),.cin(fca[953]),.sum(z[57]),.carry(fca[954]));
FA FA955 (.a(fsu[903]),.b(fca[902]),.cin(fca[954]),.sum(z[58]),.carry(fca[955]));
FA FA956 (.a(fsu[904]),.b(fca[903]),.cin(fca[955]),.sum(z[59]),.carry(fca[956]));
FA FA957 (.a(fsu[905]),.b(fca[904]),.cin(fca[956]),.sum(z[60]),.carry(fca[957]));
FA FA958 (.a(fsu[906]),.b(fca[905]),.cin(fca[957]),.sum(z[61]),.carry(fca[958]));
FA FA959 (.a(hsu[156]),.b(fca[906]),.cin(fca[958]),.sum(z[62]),.carry(fca[959]));
HA HA158 (.a(hca[156]),.b(fca[959]),.sum_h(z[63]),.carry_h(z[64]));
endmodule
