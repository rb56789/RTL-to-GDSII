`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/12/2024 02:25:41 PM
// Design Name: 
// Module Name: DA_16
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module half_adder (
    input a,b,
    output sum,carry
);

xor o1(sum,a,b);

and a1(carry,a,b);
    
endmodule

module full_adder (
    input a,b,c,
    output sum,carry
);

wire [2:0] y;

xor o1(y[0],a,b);
xor o2(sum,y[0],c);

and a1(y[1],a,b);
and a2(y[2],c,y[0]);

or o3(carry,y[1],y[2]);
    
endmodule


module com4_2 (
    input a,b,c,d,cin,
    output sum,cout,carry
);

wire [7:0] y;

xor o1(y[0],a,b);
xor o2(y[1],c,y[0]);
xor o3(y[2],d,y[1]);
xor o4(sum,cin,y[2]);

and a1(y[3],a,b);
and a2(y[4],c,y[0]);
or a3(cout,y[3],y[4]);

and a4(y[5],y[1],d);
and a5(y[6],y[2],cin);

or a6(carry,y[5],y[6]);

endmodule


module com3_2 (
    input a,b,c,cin,
    output sum,cout,carry
);

wire [6:0] y;

xor o1(y[0],a,b);
xor o2(y[1],c,y[0]);
xor o3(sum,cin,y[1]);


and a1(y[2],a,b);
and a2(y[3],c,y[0]);
or a3(cout,y[2],y[3]);

and a4(carry,y[1],cin);
    
endmodule


module DA_16 (
    input [15:0] a,b,
    output [31:0] z
);

wire [200:0] s,co,c;

wire [0:15] p[0:15];

genvar g,k;

generate
    for (g = 0; g<16; g=g+1) begin
        for (k = 0; k<16; k=k+1) begin
            and a1(p[g][k],a[k],b[g]);
        end
    end
endgenerate

//code writing 
half_adder a1(p[0][7],p[1][6],s[0],co[0]);


com3_2 a2(p[0][8],p[1][7],p[2][6],co[0],      s[1],co[1],c[0]);


com4_2 a3(p[0][9],p[1][8],p[2][7],p[3][6],co[1],     s[2],co[2],c[1]);
half_adder a4(p[4][5],p[5][4],                       s[3],co[3]);


com4_2 a5(p[0][10],p[1][9],p[2][8],p[3][7],co[2],      s[4],co[4],c[2]);
com3_2 a6(p[4][6],p[5][5],p[6][4],co[3],               s[5],co[5],c[3]);


com4_2 a7(p[0][11],p[1][10],p[2][9],p[3][8],co[4],      s[6],co[6],c[4]);
com4_2 a8(p[4][7],p[5][6],p[6][5],p[7][4],co[5],         s[7],co[7],c[5]);
half_adder a9(p[8][3],p[9][2],                           s[8],co[8]);


com4_2 a10(p[0][12],p[1][11],p[2][10],p[3][9],co[6],     s[9],co[9],c[6]);
com4_2 a11(p[4][8],p[5][7],p[6][6],p[7][5],co[7],         s[10],co[10],c[7]);
com3_2 a12(p[8][4],p[9][3],p[10][2],co[8],                s[11],co[11],c[8]);


com4_2 a13(p[0][13],p[1][12],p[2][11],p[3][10],co[9],      s[12],co[12],c[9]);
com4_2 a14(p[4][9],p[5][8],p[6][7],p[7][6],co[10],         s[13],co[13],c[10]);
com4_2 a15(p[8][5],p[9][4],p[10][3],p[11][2],co[11],       s[14],co[14],c[11]);
half_adder a16(p[12][1],p[13][0],                          s[15],co[15]);


com4_2 a17(p[0][14],p[1][13],p[2][12],p[3][11],co[12],      s[16],co[16],c[12]);
com4_2 a18(p[4][10],p[5][9],p[6][8],p[7][7],co[13],         s[17],co[17],c[13]);
com4_2 a19(p[8][6],p[9][5],p[10][4],p[11][3],co[14],        s[18],co[18],c[14]);
com3_2 a20(p[12][2],p[13][1],p[14][0],co[15],                s[19],co[19],c[15]);


com4_2 a21(p[0][15],p[1][14],p[2][13],p[3][12],co[16],       s[20],co[20],c[16]);
com4_2 a22(p[4][11],p[5][10],p[6][9],p[7][8],co[17],          s[21],co[21],c[17]);
com4_2 a23(p[8][7],p[9][6],p[10][5],p[11][4],co[18],         s[22],co[22],c[18]);
com4_2 a24(p[12][3],p[13][2],p[14][1],p[15][0],co[19],        s[23],co[23],co[24]);




com4_2 a25(p[1][15],p[2][14],p[3][13],p[4][12],co[20],        s[24],co[25],c[19]);
com4_2 a26(p[5][11],p[6][10],p[7][9],p[8][8],co[21],          s[25],co[26],c[20]);
com4_2 a27(p[9][7],p[10][6],p[11][5],p[12][4],co[22],         s[26],co[27],c[21]);
com4_2 a28(p[13][3],p[14][2],p[15][1],co[23],co[24],          s[27],co[28],co[29]);

com4_2 a29(p[2][15],p[3][14],p[4][13],p[5][12],co[25],         s[28],co[30],c[22]);
com4_2 a30(p[6][11],p[7][10],p[8][9],p[9][8],co[26],            s[29],co[31],c[23]);
com4_2 a31(p[10][7],p[11][6],p[12][5],p[13][4],co[27],          s[30],co[32],c[24]);
com3_2 a32(p[14][3],p[15][2],co[28],co[29],                     s[31],co[33],co[34]);

com4_2 a33(p[3][15],p[4][14],p[5][13],p[6][12],co[30],          s[32],co[35],c[25]);
com4_2 a34(p[7][11],p[8][10],p[9][9],p[10][8],co[31],           s[33],co[36],c[26]);
com4_2 a35(p[11][7],p[12][6],p[13][5],p[14][4],co[32],           s[34],co[37],c[27]);
full_adder a36(p[15][3],co[33],co[34],                          s[35],c[28]);

com4_2 a37(p[4][15],p[5][14],p[6][13],p[7][12],co[35],          s[36],co[38],c[29]);
com4_2 a38(p[8][11],p[9][10],p[10][9],p[11][8],co[36],          s[37],co[39],c[30]);
com4_2 a39(p[12][7],p[13][6],p[14][5],p[15][4],co[37],          s[38],co[40],c[31]);

com4_2 a40(p[5][15],p[6][14],p[7][13],p[8][12],co[38],          s[39],co[41],c[32]);
com3_2 a41(p[9][11],p[10][10],p[11][9],co[39],                  s[40],co[42],c[33]);
com3_2 a42(p[12][8],p[13][7],p[14][6],co[40],                   s[41],co[43],c[34]);

com3_2 a43(p[6][15],p[7][14],p[8][13],co[41],                   s[42],co[44],c[35]);
com3_2 a44(p[9][12],p[10][11],p[11][10],co[42],                  s[43],co[45],c[36]);
com3_2 a45(p[12][9],p[13][8],p[14][7],co[43],                    s[44],co[46],c[37]);

com3_2 a46(p[7][15],p[8][14],p[9][13],co[44],                    s[45],co[47],c[38]);
com3_2 a47(p[10][12],p[11][11],p[12][10],co[45],                 s[46],co[48],c[39]);
full_adder a48(p[13][9],p[14][8],co[46],                         s[47],c[40]);

com3_2 a49 (p[8][15],p[9][14],p[10][13],co[47],                  s[48],co[49],c[41]);
full_adder a50(p[11][12],p[12][11],co[48],                        s[49],c[42]);
half_adder a51(p[13][10],p[14][9],                                s[50],c[43]);


full_adder a52(p[9][15],p[10][14],co[49],                         s[51],c[44]);
half_adder a53(p[11][13],p[12][12],                               s[52],c[45]);
half_adder a54(p[13][11],p[14][10],                                s[53],c[46]);

half_adder a55(p[10][15],p[11][14],                               s[54],c[47]);
half_adder a56(p[12][13],p[13][12],                               s[55],c[48]);




//stage 2:
half_adder b1(p[0][2],p[1][1],                                    s[56],co[50]);


com3_2      b2(p[0][3],p[1][2],p[2][1],co[50],                    s[57],co[51],c[49]);


com4_2      b3(p[0][4],p[1][3],p[2][2],p[3][1],co[51],            s[58],co[52],c[50]);

com4_2      b4(p[0][5],p[1][4],p[2][3],p[3][2],co[52],            s[59],co[53],c[51]);
half_adder  b5(p[4][1],p[5][0],                                   s[60],co[54]);

com4_2      b6(p[0][6],p[1][5],p[2][4],p[3][3],co[53],            s[61],co[55],c[52]);
com3_2      b7(p[4][2],p[5][1],p[6][0],co[54],                    s[62],co[56],c[53]);

com4_2      b8(s[0],p[2][5],p[3][4],p[4][3],co[55],               s[63],co[57],c[54]);
com3_2      b9(p[5][2],p[6][1],p[7][0],co[56],                    s[64],co[58],c[55]);

com4_2      b10(s[1],p[3][5],p[4][4],p[5][3],co[57],              s[65],co[59],c[56]);
com3_2     b11(p[6][2],p[7][1],p[8][0],co[58],                    s[66],co[60],c[57]);

com4_2     b12(s[2],s[3],c[0],p[6][3],co[59],                 s[67],co[61],c[58]);
com3_2     b13(p[7][2],p[8][1],p[9][0],co[60],                s[68],co[62],c[59]);

com4_2     b14(s[4],s[5],c[1],p[7][3],co[61],                 s[69],co[63],c[60]);
com3_2     b15(p[8][2],p[9][1],p[10][0],co[62],                s[70],co[64],c[61]);

com4_2     b16(s[6],s[7],s[8],c[2],co[63],                   s[71],co[65],c[62]);
com3_2     b17(c[3],p[10][1],p[11][0],co[64],                s[72],co[66],c[63]);

com4_2     b18(s[9],s[10],s[11],c[4],co[65],                 s[73],co[67],c[64]);
com3_2     b19(c[5],p[11][1],p[12][0],co[66],                s[74],co[68],c[65]);

com4_2     b20(s[12],s[13],s[14],s[15],co[67],               s[75],co[69],c[66]);
com3_2     b21(c[6],c[7],c[8],co[68],                        s[76],co[70],c[67]);

com4_2     b22(s[16],s[17],s[18],s[19],co[69],               s[77],co[71],c[68]);
com3_2     b23(c[9],c[10],c[11],co[70],                      s[78],co[72],c[69]);

com4_2     b24(s[20],s[21],s[22],s[23],co[71],               s[79],co[73],c[70]);
com4_2     b25(c[12],c[13],c[14],c[15],co[72],               s[80],co[74],c[71]);

com4_2     b26(s[24],s[25],s[26],s[27],co[73],               s[81],co[75],c[72]);
com3_2     b27(c[16],c[17],c[18],co[74],                     s[82],co[76],c[73]);

com4_2     b28(s[28],s[29],s[30],s[31],co[75],               s[83],co[77],c[74]);
com3_2     b29(c[19],c[20],c[21],co[76],                     s[84],co[78],c[75]);

com4_2     b30(s[32],s[33],s[34],s[35],co[77],               s[85],co[79],c[76]);
com3_2     b31(c[22],c[23],c[24],co[78],                     s[86],co[80],c[77]);

com4_2     b32(s[36],s[37],s[38],c[25],co[79],               s[87],co[81],c[78]);
com3_2     b33(c[26],c[27],c[28],co[80],                     s[88],co[82],c[79]);

com4_2     b34(s[39],s[40],s[41],p[15][5],co[81],            s[89],co[83],c[80]);
com3_2     b35(c[29],c[30],c[31],co[82],                     s[90],co[84],c[81]);

com4_2    b36(s[42],s[43],s[44],p[15][6],co[83],             s[91],co[85],c[82]);
com3_2    b37(c[32],c[33],c[34],co[84],                      s[92],co[86],c[83]);

com4_2    b38(s[45],s[46],s[47],p[15][7],co[85],             s[93],co[87],c[84]);
com3_2    b39(c[35],c[36],c[37],co[86],                      s[94],co[88],c[85]);

com4_2    b40(s[48],s[49],s[50],p[15][8],co[87],             s[95],co[89],c[86]);
com3_2    b41(c[38],c[39],c[40],co[88],                      s[96],co[90],c[87]);

com4_2    b42(s[51],s[52],s[53],p[15][9],co[89],             s[97],co[91],c[88]);
com3_2    b43(c[41],c[42],c[43],co[90],                      s[98],co[92],c[89]);

com4_2    b44(s[54],s[55],p[14][11],p[15][10],co[91],        s[99],co[93],c[90]);
com3_2    b45(c[44],c[45],c[46],co[92],                      s[100],co[94],c[91]);

com4_2    b46(p[11][15],p[12][14],p[13][13],p[14][12],co[93], s[101],co[95],c[92]);
com3_2    b47(p[15][11],c[47],c[48],co[94],                   s[102],co[96],c[93]);

full_adder b48(p[12][15],p[13][14],co[95],                    s[103],co[97]);
full_adder b49(p[14][13],p[15][12],co[96],                    s[104],co[98]);

half_adder b50(p[13][15],co[97],                              s[105],c[94]);
full_adder b51(p[14][14],p[15][13],co[98],                    s[106],co[99]);

full_adder b52(p[14][15],p[15][14],co[99],                    s[107],c[95]);


//stage 3:

assign z[0]=p[0][0];
half_adder c1(p[0][1],p[1][0],           z[1],co[100]);
full_adder c2(s[56],p[2][0],co[100],     z[2],co[101]);
full_adder c3(s[57],p[3][0],co[101],     z[3],co[102]);
com3_2 c4(s[58],c[49],p[4][0],co[102],   z[4],co[103],c[96]);
com3_2 c5(s[59],s[60]      ,c[50],co[103],      s[108],co[104],c[97]);
com3_2 c6(s[61],s[62]      ,c[51],  co[104],      s[109],co[105],c[98]);
com4_2 c7(s[63],s[64],c[52],c[53],co[105],s[110],co[106],c[99]);
com4_2 c8(s[65],s[66],c[54],c[55],co[106],s[111],co[107],c[100]);
com4_2 c9(s[67],s[68],c[56],c[57],co[107],s[112],co[108],c[101]);
com4_2 c10(s[69],s[70],c[58],c[59],co[108],s[113],co[109],c[102]);
com4_2 c11(s[71],s[72],c[60],c[61],co[109],s[114],co[110],c[103]);
com4_2 c12(s[73],s[74],c[62],c[63],co[110],s[115],co[111],c[104]);
com4_2 c13(s[75],s[76],c[64],c[65],co[111],s[116],co[112],c[105]);
com4_2 c14(s[77],s[78],c[66],c[67],co[112],s[117],co[113],c[106]);
com4_2 c15(s[79],s[80],c[68],c[69],co[113],s[118],co[114],c[107]);
com4_2 c16(s[81],s[82],c[70],c[71],co[114],s[119],co[115],c[108]);
com4_2 c17(s[83],s[84],c[72],c[73],co[115],s[120],co[116],c[109]);
com4_2 c18(s[85],s[86],c[74],c[75],co[116],s[121],co[117],c[110]);
com4_2 c19(s[87],s[88],c[76],c[77],co[117],s[122],co[118],c[111]);
com4_2 c20(s[89],s[90],c[78],c[79],co[118],s[123],co[119],c[112]);
com4_2 c21(s[91],s[92],c[80],c[81],co[119],s[124],co[120],c[113]);
com4_2 c22(s[93],s[94],c[82],c[83],co[120],s[125],co[121],c[114]);
com4_2 c23(s[95],s[96],c[84],c[85],co[121],s[126],co[122],c[115]);
com4_2 c24(s[97],s[98],c[86],c[87],co[122],s[127],co[123],c[116]);
com4_2 c25(s[99],s[100],c[88],c[89],co[123],s[128],co[124],c[117]);
com4_2 c26(s[101],s[102],c[90],c[91],co[124],s[129],co[125],c[118]);
com4_2 c27(s[103],s[104],c[92],c[93],co[125],s[130],co[126],c[119]);

full_adder c28(s[105],s[106],co[126],        s[131],c[120]);
full_adder d1(s[107],c[94],c[120],           s[132],c[121]);
full_adder d2(p[15][15],c[95],c[121],        s[133],c[122]);



half_adder e29(s[108],c[96],         z[5],co[127]);
full_adder c29(s[109],c[97],co[127],        z[6],co[128]);
full_adder c30(s[110],co[128],c[98 ], z[7], co[129]);
full_adder c31(s[111],co[129],c[99 ], z[8], co[130]);
full_adder c32(s[112],co[130],c[100], z[9], co[131]);
full_adder c33(s[113],co[131],c[101],z[10],co[132]);
full_adder c34(s[114],co[132],c[102],z[11],co[133]);
full_adder c35(s[115],co[133],c[103],z[12],co[134]);
full_adder c36(s[116],co[134],c[104],z[13],co[135]);
full_adder c37(s[117],co[135],c[105],z[14],co[136]);
full_adder c38(s[118],co[136],c[106],z[15],co[137]);
full_adder c39(s[119],co[137],c[107],z[16],co[138]);
full_adder c40(s[120],co[138],c[108],z[17],co[139]);
full_adder c41(s[121],co[139],c[109],z[18],co[140]);
full_adder c42(s[122],co[140],c[110],z[19],co[141]);
full_adder c43(s[123],co[141],c[111],z[20],co[142]);
full_adder c44(s[124],co[142],c[112],z[21],co[143]);
full_adder c45(s[125],co[143],c[113],z[22],co[144]);
full_adder c46(s[126],co[144],c[114],z[23],co[145]);
full_adder c47(s[127],co[145],c[115],z[24],co[146]);
full_adder c48(s[128],co[146],c[116],z[25],co[147]);
full_adder c49(s[129],co[147],c[117],z[26],co[148]);
full_adder c50(s[130],co[148],c[118],z[27],co[149]);
full_adder c51(s[131],co[149],c[119],z[28],co[150]);
half_adder c52(s[132],co[150],       z[29],co[151]);
half_adder c53(s[133],co[151],       z[30],co[152]);
half_adder c54(c[122],co[152],       z[31],co[153]);





endmodule