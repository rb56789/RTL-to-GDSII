`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/20/2024 04:54:22 PM
// Design Name: 
// Module Name: DA_32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module com3_2 (
    input a,b,c,cin,
    output sum,cout,carry
);

wire [6:0] y;

xor o1(y[0],a,b);
xor o2(y[1],c,y[0]);
xor o3(sum,cin,y[1]);


and a1(y[2],a,b);
and a2(y[3],c,y[0]);
or a3(cout,y[2],y[3]);

and a4(carry,y[1],cin);
    
endmodule

module com4_2 (
    input a,b,c,d,cin,
    output sum,cout,carry
);

wire [7:0] y;

xor o1(y[0],a,b);
xor o2(y[1],c,y[0]);
xor o3(y[2],d,y[1]);
xor o4(sum,cin,y[2]);

and a1(y[3],a,b);
and a2(y[4],c,y[0]);
or a3(cout,y[3],y[4]);

and a4(y[5],y[1],d);
and a5(y[6],y[2],cin);

or a6(carry,y[5],y[6]);

endmodule

module full_adder (
    input a,b,c,
    output sum,carry
);

wire [2:0] y;

xor o1(y[0],a,b);
xor o2(sum,y[0],c);

and a1(y[1],a,b);
and a2(y[2],c,y[0]);

or o3(carry,y[1],y[2]);
    
endmodule

module half_adder (
    input a,b,
    output sum,carry
);

xor o1(sum,a,b);

and a1(carry,a,b);
    
endmodule

module DA_32 (
    input [31:0] a,b,
    output [63:0] z
);

wire [600:0] s,co,c;

wire [0:31] p[0:31];

genvar g,k;

generate
    for (g = 0; g<32; g=g+1) begin
        for (k = 0; k<32; k=k+1) begin
            and a1(p[g][k],a[k],b[g]);
        end
    end
endgenerate

//code writing 


half_adder a1(p[0][8],p[1][7],s[0],co[0]);


com3_2     a2(p[0][9],p[1][8],p[2][7],co[0], s[1],co[1],c[0]);


com4_2     a3(p[0][10],p[1][9],p[2][8],p[3][7],co[1],s[2],co[2],c[1]);

com4_2     a4(p[0][11],p[1][10],p[2][9],p[3][8],co[2],s[3],co[3],c[2]);
half_adder a5(p[4][7],p[5][6],                        s[4],co[4]);

com4_2     a6(p[0][12],p[1][11],p[2][10],p[3][9],co[3],s[5],co[5],c[3]);
com3_2     a7(p[4][8],p[5][7],p[6][6],co[4],           s[6],co[6],c[4]);

com4_2     a8(p[0][13],p[1][12],p[2][11],p[3][10],co[5],s[7],co[7],c[5]);
com4_2     a9(p[4][9],p[5][8],p[6][7],p[7][6],co[6],    s[8],co[8],c[6]);

com4_2     a10(p[0][14],p[1][13],p[2][12],p[3][11],co[7],s[9],co[9],c[7]);
com4_2     a11(p[4][10],p[5][9],p[6][8],p[7][7],co[8],   s[10],co[10],c[8]);
half_adder a12(p[8][6],p[9][5],                          s[11],co[11]);


com4_2    a13(p[0][15],p[1][14],p[2][13],p[3][12],co[9], s[12],co[12],c[9]);
com4_2    a14(p[4][11],p[5][10],p[6][9],p[7][8],co[10],  s[13],co[13],c[10]);
com3_2    a15(p[8][7],p[9][6],p[10][5],co[11],           s[14],co[14],c[11]);

com4_2    a16(p[0][16],p[1][15],p[2][14],p[3][13],co[12], s[15],co[15],c[12]);
com4_2    a17(p[4][12],p[5][11],p[6][10],p[7][9],co[13],  s[16],co[16],c[13]);
com4_2    a18(p[8][8],p[9][7],p[10][6],p[11][5],co[14],   s[17],co[17],c[14]);

com4_2    a19(p[0][17],p[1][16],p[2][15],p[3][14],co[15], s[18],co[18],c[15]);
com4_2    a20(p[4][13],p[5][12],p[6][11],p[7][10],co[16], s[19],co[19],c[16]);
com4_2    a21(p[8][9],p[9][8],p[10][7],p[11][6],co[17],   s[20],co[20],c[17]);
half_adder a22(p[12][5],p[13][4],                         s[21],co[21]);


com4_2    a23(p[0][18],p[1][17],p[2][16],p[3][15],co[18], s[22],co[22],c[18]);
com4_2    a24(p[4][14],p[5][13],p[6][12],p[7][11],co[19], s[23],co[23],c[19]);
com4_2    a25(p[8][10],p[9][9],p[10][8],p[11][7],co[20],  s[24],co[24],c[20]);
com3_2    a26(p[12][6],p[13][5],p[14][4],      co[21],     s[25],co[25],c[21]);


com4_2    a27(p[0][19],p[1][18],p[2][17],p[3][16],co[22],  s[26],co[26],c[22]);
com4_2    a28(p[4][15],p[5][14],p[6][13],p[7][12],co[23],  s[27],co[27],c[23]);
com4_2    a29(p[8][11],p[9][10],p[10][9],p[11][8],co[24],  s[28],co[28],c[24]);
com4_2    a30(p[12][7],p[13][6],p[14][5],p[15][4],co[25],  s[29],co[29],c[25]);


com4_2   a31(p[0][20],p[1][19],p[2][18],p[3][17],co[26],    s[30],co[30],c[26]);
com4_2   a32(p[4][16],p[5][15],p[6][14],p[7][13],co[27],    s[31],co[31],c[27]);
com4_2   a33(p[8][12],p[9][11],p[10][10],p[11][9],co[28],   s[32],co[32],c[28]);
com4_2   a34(p[12][8],p[13][7],p[14][6],p[15][5],co[29],    s[33],co[33],c[29]);
half_adder a35(p[16][4],p[17][3],                           s[34],co[34]);

com4_2 a36(p[0][21],p[1][20],p[2][19],p[3][18],co[30],      s[35],co[35],c[30]);
com4_2 a37(p[4][17],p[5][16],p[6][15],p[7][14],co[31],      s[36],co[36],c[31]);
com4_2 a38(p[8][13],p[9][12],p[10][11],p[11][10],co[32],    s[37],co[37],c[32]);
com4_2 a39(p[12][9],p[13][8],p[14][7],p[15][6],co[33],      s[38],co[38],c[33]);
com3_2 a40(p[16][5],p[17][4],p[18][3],co[34],               s[39],co[39],c[34]);

com4_2 a41(p[0][22],p[1][21],p[2][20],p[3][19],co[35],      s[40],co[40],c[35]);
com4_2 a42(p[4][18],p[5][17],p[6][16],p[7][15],co[36],      s[41],co[41],c[36]);
com4_2 a43(p[8][14],p[9][13],p[10][12],p[11][11],co[37],    s[42],co[42],c[37]);
com4_2 a44(p[12][10],p[13][9],p[14][8],p[15][7],co[38],     s[43],co[43],c[38]);
com4_2 a45(p[16][6],p[17][5],p[18][4],p[19][3],co[39],      s[44],co[44],c[39]);

com4_2 a46(p[0][23],p[1][22],p[2][21],p[3][20],co[40],      s[45],co[45],c[40]);
com4_2 a47(p[4][19],p[5][18],p[6][17],p[7][16],co[41],      s[46],co[46],c[41]);
com4_2 a48(p[8][15],p[9][14],p[10][13],p[11][12],co[42],    s[47],co[47],c[42]);
com4_2 a49(p[12][11],p[13][10],p[14][9],p[15][8],co[43],     s[48],co[48],c[43]);
com4_2 a50(p[16][7],p[17][6],p[18][5],p[19][4],co[44],      s[49],co[49],c[44]);
half_adder a51(p[20][3],p[21][2],                            s[50],co[50]);

com4_2 a52(p[0][24],p[1][23],p[2][22],p[3][21],co[45],      s[51],co[51],c[45]);
com4_2 a53(p[4][20],p[5][19],p[6][18],p[7][17],co[46],      s[52],co[52],c[46]);
com4_2 a54(p[8][16],p[9][15],p[10][14],p[11][13],co[47],    s[53],co[53],c[47]);
com4_2 a55(p[12][12],p[13][11],p[14][10],p[15][9],co[48],     s[54],co[54],c[48]);
com4_2 a56(p[16][8],p[17][7],p[18][6],p[19][5],co[49],      s[55],co[55],c[49]);
com3_2 a57(p[20][4],p[21][3],p[22][2],co[50],               s[56],co[56],c[50]);

com4_2 a58(p[0][25],p[1][24],p[2][23],p[3][22],co[51],      s[57],co[57],c[51]);
com4_2 a59(p[4][21],p[5][20],p[6][19],p[7][18],co[52],      s[58],co[58],c[52]);
com4_2 a60(p[8][17],p[9][16],p[10][15],p[11][14],co[53],    s[59],co[59],c[53]);
com4_2 a61(p[12][13],p[13][12],p[14][11],p[15][10],co[54],  s[60],co[60],c[54]);
com4_2 a62(p[16][9],p[17][8],p[18][7],p[19][6],co[55],      s[61],co[61],c[55]);
com4_2 a63(p[20][5],p[21][4],p[22][3],p[23][2],co[56],      s[62],co[62],c[56]);

com4_2 a64(p[0][26],p[1][25],p[2][24],p[3][23],co[57],      s[63],co[63],c[57]);
com4_2 a65(p[4][22],p[5][21],p[6][20],p[7][19],co[58],      s[64],co[64],c[58]);
com4_2 a66(p[8][18],p[9][17],p[10][16],p[11][15],co[59],    s[65],co[65],c[59]);
com4_2 a67(p[12][14],p[13][13],p[14][12],p[15][11],co[60],  s[66],co[66],c[60]);
com4_2 a68(p[16][10],p[17][9],p[18][8],p[19][7],co[61],      s[67],co[67],c[61]);
com4_2 ab67(p[20][6],p[21][5],p[22][4],p[23][3],co[62],      s[68],co[68],c[62]);
half_adder ab68(p[24][2],p[25][1],                           s[69],co[69]);

com4_2 a69(p[0][27],p[1][26],p[2][25],p[3][24],co[63],      s[70],co[70],c[63]);
com4_2 a70(p[4][23],p[5][22],p[6][21],p[7][20],co[64],      s[71],co[71],c[64]);
com4_2 a71(p[8][19],p[9][18],p[10][17],p[11][16],co[65],    s[72],co[72],c[65]);
com4_2 a72(p[12][15],p[13][14],p[14][13],p[15][12],co[66],  s[73],co[73],c[66]);
com4_2 a73(p[16][11],p[17][10],p[18][9],p[19][8],co[67],    s[74],co[74],c[67]);
com4_2 a74(p[20][7],p[21][6],p[22][5],p[23][4],co[68],      s[75],co[75],c[68]);
com3_2 a75(p[24][3],p[25][2],p[26][1],co[69],               s[76],co[76],c[69]);

com4_2 a76(p[0][28],p[1][27],p[2][26],p[3][25],co[70],      s[77],co[77],c[70]);
com4_2 a77(p[4][24],p[5][23],p[6][22],p[7][21],co[71],      s[78],co[78],c[71]);
com4_2 a78(p[8][20],p[9][19],p[10][18],p[11][17],co[72],   s[79],co[79],c[72]);
com4_2 a79(p[12][16],p[13][15],p[14][14],p[15][13],co[73],  s[80],co[80],c[73]);
com4_2 a80(p[16][12],p[17][11],p[18][10],p[19][9],co[74],   s[81],co[81],c[74]);
com4_2 a81(p[20][8],p[21][7],p[22][6],p[23][5],co[75],      s[82],co[82],c[75]);
com4_2 a82(p[24][4],p[25][3],p[26][2],p[27][1],co[76],      s[83],co[83],c[76]);

com4_2 a83(p[0][29],p[1][28],p[2][27],p[3][26],co[77],      s[84],co[84],c[77]);
com4_2 a84(p[4][25],p[5][24],p[6][23],p[7][22],co[78],      s[85],co[85],c[78]);
com4_2 a85(p[8][21],p[9][20],p[10][19],p[11][18],co[79],   s[86],co[86],c[79]);
com4_2 a86(p[12][17],p[13][16],p[14][15],p[15][14],co[80],  s[87],co[87],c[80]);
com4_2 a87(p[16][13],p[17][12],p[18][11],p[19][10],co[81],   s[88],co[88],c[81]);
com4_2 a88(p[20][9],p[21][8],p[22][7],p[23][6],co[82],      s[89],co[89],c[82]);
com4_2 a89(p[24][5],p[25][4],p[26][3],p[27][2],co[83],      s[90],co[90],c[83]);
half_adder a90(p[28][1],p[29][0],                           s[91],co[91]);

com4_2 a91(p[0][30],p[1][29],p[2][28],p[3][27],co[84],      s[92],co[92],c[85]);
com4_2 a92(p[4][26],p[5][25],p[6][24],p[7][23],co[85],      s[93],co[93],c[86]);
com4_2 a93(p[8][22],p[9][21],p[10][20],p[11][19],co[86],   s[94],co[94],c[87]);
com4_2 a94(p[12][18],p[13][17],p[14][16],p[15][15],co[87],  s[95],co[95],c[88]);
com4_2 a95(p[16][14],p[17][13],p[18][12],p[19][11],co[88],   s[96],co[96],c[89]);
com4_2 a96(p[20][10],p[21][9],p[22][8],p[23][7],co[89],      s[97],co[97],c[90]);
com4_2 a97(p[24][6],p[25][5],p[26][4],p[27][3],co[90],      s[98],co[98],c[91]);
com3_2 a98(p[28][2],p[29][1],p[30][0],co[91],               s[99],co[99],c[92]);

com4_2 a99(p[0][31],p[1][30],p[2][29],p[3][28],co[92],      s[100],co[100],c[93]);
com4_2 a100(p[4][27],p[5][26],p[6][25],p[7][24],co[93],      s[101],co[101],c[94]);
com4_2 a101(p[8][23],p[9][22],p[10][21],p[11][20],co[94],   s[102],co[102],c[95]);
com4_2 a102(p[12][19],p[13][18],p[14][17],p[15][16],co[95],  s[103],co[103],c[96]);
com4_2 a103(p[16][15],p[17][14],p[18][13],p[19][12],co[96],   s[104],co[104],c[97]);
com4_2 a104(p[20][11],p[21][10],p[22][9],p[23][8],co[97],      s[105],co[105],c[98]);
com4_2 a105(p[24][7],p[25][6],p[26][5],p[27][4],co[98],      s[106],co[106],c[99]);
com4_2 a106(p[28][3],p[29][2],p[30][1],p[31][0],co[99],      s[107],co[107],co[108]);

com4_2 a107(p[1][31],p[2][30],p[3][29],p[4][28],co[100],     s[108],co[109],c[100]);
com4_2 a108(p[5][27],p[6][26],p[7][25],p[8][24],co[101],     s[109],co[110],c[101]);
com4_2 a109(p[9][23],p[10][22],p[11][21],p[12][20],co[102],  s[110],co[111],c[102]);
com4_2 a110(p[13][19],p[14][18],p[15][17],p[16][16],co[103], s[111],co[112],c[103]);
com4_2 a111(p[17][15],p[18][14],p[19][13],p[20][12],co[104], s[112],co[113],c[104]);
com4_2 a112(p[21][11],p[22][10],p[23][9],p[24][8],co[105],   s[113],co[114],c[105]);
com4_2 a113(p[25][7],p[26][6],p[27][5],p[28][4],co[106],     s[114],co[115],c[106]);
com4_2 a114(p[29][3],p[30][2],p[31][1],co[107],co[108],      s[115],co[116],co[117]);

com4_2 a115(p[2][31],p[3][30],p[4][29],p[5][28],co[109],     s[116],co[118],c[107]);
com4_2 a116(p[6][27],p[7][26],p[8][25],p[9][24],co[110],     s[117],co[119],c[108]);
com4_2 a117(p[10][23],p[11][22],p[12][21],p[13][20],co[111],  s[118],co[120],c[109]);
com4_2 a118(p[14][19],p[15][18],p[16][17],p[17][16],co[112], s[119],co[121],c[110]);
com4_2 a119(p[18][15],p[19][14],p[20][13],p[21][12],co[113], s[120],co[122],c[111]);
com4_2 a120(p[22][11],p[23][10],p[24][9],p[25][8],co[114],   s[121],co[123],c[112]);
com4_2 a121(p[26][7],p[27][6],p[28][5],p[29][4],co[115],     s[122],co[124],c[113]);
com3_2 a122(p[30][3],p[31][2],co[116],co[117],               s[123],co[125],co[126]);

com4_2 a123(p[3][31],p[4][30],p[5][29],p[6][28],co[118],     s[124],co[127],c[114]);
com4_2 a124(p[7][27],p[8][26],p[9][25],p[10][24],co[119],     s[125],co[128],c[115]);
com4_2 a125(p[11][23],p[12][22],p[13][21],p[14][20],co[120],  s[126],co[129],c[116]);
com4_2 a126(p[15][19],p[16][18],p[17][17],p[18][16],co[121], s[127],co[130],c[117]);
com4_2 a127(p[19][15],p[20][14],p[21][13],p[22][12],co[122], s[128],co[131],c[118]);
com4_2 a128(p[23][11],p[24][10],p[25][9],p[26][8],co[123],   s[129],co[132],c[119]);
com4_2 a129(p[27][7],p[28][6],p[29][5],p[30][4],co[124],     s[130],co[133],c[120]);
full_adder a130(p[31][3],co[125],co[126],                    s[131],        c[121]);

com4_2 a131(p[4][31],p[5][30],p[6][29],p[7][28],co[127],     s[132],co[134],c[122]);
com4_2 a132(p[8][27],p[9][26],p[10][25],p[11][24],co[128],     s[133],co[135],c[123]);
com4_2 a133(p[12][23],p[13][22],p[14][21],p[15][20],co[129],  s[134],co[136],c[124]);
com4_2 a134(p[16][19],p[17][18],p[18][17],p[19][16],co[130], s[135],co[137],c[125]);
com4_2 a135(p[20][15],p[21][14],p[22][13],p[23][12],co[131], s[136],co[138],c[126]);
com4_2 a136(p[24][11],p[25][10],p[26][9],p[27][8],co[132],   s[137],co[139],c[127]);
com3_2 a137(p[28][7],p[29][6],p[30][5],co[133],              s[138],co[140],c[128]);

com4_2 a138(p[5][31],p[6][30],p[7][29],p[8][28],co[134],     s[139],co[141],c[129]);
com4_2 a139(p[9][27],p[10][26],p[11][25],p[12][24],co[135],     s[140],co[142],c[130]);
com4_2 a140(p[13][23],p[14][22],p[15][21],p[16][20],co[136],  s[141],co[143],c[131]);
com4_2 a141(p[17][19],p[18][18],p[19][17],p[20][16],co[137], s[142],co[144],c[132]);
com4_2 a142(p[21][15],p[22][14],p[23][13],p[24][12],co[138], s[143],co[145],c[133]);
com4_2 a143(p[25][11],p[26][10],p[27][9],p[28][8],co[139],   s[144],co[146],c[134]);
full_adder a144(p[29][7],p[30][6],co[140],                   s[145],        c[135]);

com4_2 a145(p[6][31],p[7][30],p[8][29],p[9][28],co[141],     s[146],co[147],c[136]);
com4_2 a146(p[10][27],p[11][26],p[12][25],p[13][24],co[142],     s[147],co[148],c[137]);
com4_2 a147(p[14][23],p[15][22],p[16][21],p[17][20],co[143],  s[148],co[149],c[138]);
com4_2 a148(p[18][19],p[19][18],p[20][17],p[21][16],co[144], s[149],co[150],c[139]);
com4_2 a149(p[22][15],p[23][14],p[24][13],p[25][12],co[145], s[150],co[151],c[140]);
com4_2 a150(p[26][11],p[27][10],p[28][9],p[29][8],co[146],   s[151],co[152],c[141]);


com4_2 ab145(p[7][31],p[8][30],p[9][29],p[10][28],co[147],     s[152],co[153],c[142]);
com4_2 ab146(p[11][27],p[12][26],p[13][25],p[14][24],co[148],     s[153],co[154],c[143]);
com4_2 ab147(p[15][23],p[16][22],p[17][21],p[18][20],co[149],  s[154],co[155],c[144]);
com4_2 ab148(p[19][19],p[20][18],p[21][17],p[22][16],co[150], s[155],co[156],c[145]);
com4_2 ab149(p[23][15],p[24][14],p[25][13],p[26][12],co[151], s[156],co[157],c[146]);
full_adder ab150(p[27][11],p[28][10],co[152],                     s[157],        c[147]);


com4_2 a151(p[8][31],p[9][30],p[10][29],p[11][28],co[153],     s[158],co[158],c[148]);
com4_2 a152(p[12][27],p[13][26],p[14][25],p[15][24],co[154],     s[159],co[159],c[149]);
com4_2 a153(p[16][23],p[17][22],p[18][21],p[19][20],co[155],  s[160],co[160],c[150]);
com4_2 a154(p[20][19],p[21][18],p[22][17],p[23][16],co[156], s[161],co[161],c[151]);
com4_2 a155(p[24][15],p[25][14],p[26][13],p[27][12],co[157], s[162],co[162],c[152]);


com4_2 a156(p[9][31],p[10][30],p[11][29],p[12][28],co[158],     s[163],co[163],c[153]);
com4_2 a157(p[13][27],p[14][26],p[15][25],p[16][24],co[159],     s[164],co[164],c[154]);
com4_2 a158(p[17][23],p[18][22],p[19][21],p[20][20],co[160],  s[165],co[165],c[155]);
com4_2 a159(p[21][19],p[22][18],p[23][17],p[24][16],co[161], s[166],co[166],c[156]);
full_adder a160(p[25][15],p[26][14],co[162],                     s[167],        c[157]);


com4_2 a161(p[10][31],p[11][30],p[12][29],p[13][28],co[163],     s[168],co[167],c[158]);
com4_2 a162(p[14][27],p[15][26],p[16][25],p[17][24],co[164],     s[169],co[168],c[159]);
com4_2 a163(p[18][23],p[19][22],p[20][21],p[21][20],co[165],  s[170],co[169],c[160]);
com4_2 a164(p[22][19],p[23][18],p[24][17],p[25][16],co[166], s[171],co[170],c[161]);


com4_2 a165(p[11][31],p[12][30],p[13][29],p[14][28],co[167],     s[172],co[171],c[162]);
com4_2 a166(p[15][27],p[16][26],p[17][25],p[18][24],co[168],     s[173],co[172],c[163]);
com4_2 a167(p[19][23],p[20][22],p[21][21],p[22][20],co[169],     s[174],co[173],c[164]);
full_adder a168(p[23][19],p[24][18],co[170],                     s[175],        c[165]);


com4_2 a169(p[12][31],p[13][30],p[14][29],p[15][28],co[171],     s[176],co[174],c[166]);
com4_2 a170(p[16][27],p[17][26],p[18][25],p[19][24],co[172],     s[177],co[175],c[167]);
com4_2 a171(p[20][23],p[21][22],p[22][21],p[23][20],co[173],     s[178],co[176],c[168]);


com4_2 a172(p[13][31],p[14][30],p[15][29],p[16][28],co[174],     s[179],co[177],c[169]);
com4_2 a173(p[17][27],p[18][26],p[19][25],p[20][24],co[175],     s[180],co[178],c[170]);
full_adder a174(p[21][23],p[22][22],                co[176],     s[181],        c[171]);


com4_2 ab172(p[14][31],p[15][30],p[16][29],p[17][28],co[177],     s[182],co[179],c[172]);
com4_2 ab173(p[18][27],p[19][26],p[20][25],p[21][24],co[178],     s[183],co[180],c[173]);


com4_2 ab174(p[15][31],p[16][30],p[17][29],p[18][28],co[179],     s[184],co[181],c[174]);
full_adder a175(p[19][27],p[20][26]                    ,co[180],     s[185],        c[175]);


com4_2 a176(p[16][31],p[17][30],p[18][29],p[19][28],co[181],     s[186],co[182],c[176]);

full_adder a177(p[17][31],p[18][30]                    ,co[182],     s[187],c[177]);


//stage 2:
half_adder b1(p[0][2],p[1][1],s[188],co[183]);

com3_2  b2(p[0][3],p[1][2],p[2][1],co[183],   s[189],co[184],c[178]);

com4_2 b3(p[0][4],p[1][3],p[2][2],p[3][1],co[184], s[190],co[185],c[179]);

com4_2 b4(p[0][5],p[1][4],p[2][3],p[3][2],co[185], s[191],co[186],c[180]);
half_adder b5(p[4][1],p[5][0],                     s[192],co[187]);

com4_2 b6(p[0][6],p[1][5],p[2][4],p[3][3],co[186], s[193],co[188],c[181]);
com3_2 b7(p[4][2],p[5][1],p[6][0],co[187],          s[194],co[189],c[182]);

com4_2 b8(p[0][7],p[1][6],p[2][5],p[3][4],co[188],  s[195],co[190],c[183]);
com4_2 b9(p[4][3],p[5][2],p[6][1],p[7][0],co[189],  s[196],co[191],c[184]);

com4_2 b10(s[0],p[2][6],p[3][5],p[4][4],co[190],    s[197],co[192],c[185]);
com4_2 b11(p[5][3],p[6][2],p[7][1],p[8][0],co[191], s[198],co[193],c[186]);

com4_2 b12(s[1],p[3][6],p[4][5],p[5][4],co[192],     s[199],co[194],c[187]);
com4_2 b13(p[6][3],p[7][2],p[8][1],p[9][0],co[193],  s[200],co[195],c[188]);

com4_2 b14(s[2],c[0],p[4][6],p[5][5],co[194],        s[201],co[196],c[189]);
com4_2 b15(p[6][4],p[7][3],p[8][2],p[9][1],co[195],  s[202],co[197],c[190]);

com4_2 b16(s[3],s[4],c[1],p[6][5],co[196],           s[203],co[198],c[191]);
com4_2 b17(p[7][4],p[8][3],p[9][2],p[10][1],co[197], s[204],co[199],c[192]);

com4_2 b18(s[5],s[6],c[2],p[7][5],co[198],           s[205],co[200],c[193]);
com4_2 b19(p[8][4],p[9][3],p[10][2],p[11][1],co[199],s[206],co[201],c[194]);

com4_2 b20(s[7],s[8],c[3],c[4],co[200],               s[207],co[202],c[195]);
com4_2 b21(p[8][5],p[9][4],p[10][3],p[11][2],co[201], s[208],co[203],c[196]);
half_adder b22(p[12][1],p[13][0],                     s[209],co[204]);

com4_2 b23(s[9],s[10],s[11],p[10][4],co[202],          s[210],co[205],c[197]);
com4_2 b24(c[5],c[6],p[11][3],p[12][2],co[203],        s[211],co[206],c[198]);
full_adder b25(p[13][1],p[14][0],co[204],              s[212],co[207]);

com4_2 b26(s[12],s[13],s[14],p[11][4],co[205],         s[213],co[208],c[199]);
com4_2 b27(c[7],c[8],p[12][3],p[13][2],co[206],        s[214],co[209],c[200]);
full_adder b28(p[14][1],p[15][0],co[207],              s[215],co[210]);

com4_2 b29(s[15],s[16],s[17],p[12][4],co[208],         s[216],co[211],c[201]);
com4_2 b30(c[9],c[10],c[11],p[13][3],co[209],           s[217],co[212],c[202]);
com3_2 b31(p[14][2],p[15][1],p[16][0],co[210],         s[218],co[213],c[203]);

com4_2 b32(s[18],s[19],s[20],s[21],co[211],            s[219],co[214],c[204]);
com4_2 b33(c[12],c[13],c[14],p[14][3],co[212],         s[220],co[215],c[205]);
com3_2 b34(p[15][2],p[16][1],p[17][0],co[213],         s[221],co[216],c[206]);

com4_2 b35(s[22],s[23],s[24],s[25],co[214],            s[222],co[217],c[207]);
com4_2 b36(c[15],c[16],c[17],p[15][3],co[215],         s[223],co[218],c[208]);
com3_2 b37(p[16][2],p[17][1],p[18][0],co[216],         s[224],co[219],c[209]);

com4_2 b38(s[26],s[27],s[28],s[29],co[217],            s[225],co[220],c[210]);
com4_2 b39(c[18],c[19],c[20],c[21],co[218],            s[226],co[221],c[211]);
com4_2 b40(p[16][3],p[17][2],p[18][1],p[19][0],co[219], s[227],co[222],c[212]);

com4_2 b41(s[30],s[31],s[32],s[33],co[220],            s[228],co[223],c[213]);
com4_2 b42(s[34],c[22],c[23],c[24],co[221],            s[229],co[224],c[214]);
com4_2 b43(c[25],p[18][2],p[19][1],p[20][0],co[222],   s[230],co[225],c[215]);

com4_2 b44(s[35],s[36],s[37],s[38],co[223],            s[231],co[226],c[216]);
com4_2 b45(s[39],c[26],c[27],c[28],co[224],            s[232],co[227],c[217]);
com4_2 b46(c[29],p[19][2],p[20][1],p[21][0],co[225],   s[233],co[228],c[218]);

com4_2 b47(s[40],s[41],s[42],s[43],co[226],             s[234],co[229],c[219]);
com4_2 b48(s[44],c[30],c[31],c[32],co[227],             s[235],co[230],c[220]);
com4_2 b49(c[33],c[34],p[20][2],p[21][1],co[228],       s[236],co[231],c[221]);

com4_2 b50(s[45],s[46],s[47],s[48],co[229],             s[237],co[232],c[222]);
com4_2 b51(s[49],s[50],c[35],c[36],co[230],             s[238],co[233],c[223]);
com4_2 b52(c[37],c[38],c[39],p[22][1],co[231],          s[239],co[234],c[224]);

com4_2 b53(s[51],s[52],s[53],s[54],co[232],             s[240],co[235],c[225]);
com4_2 b54(s[55],s[56],c[40],c[41],co[233],             s[241],co[236],c[226]);
com4_2 b55(c[42],c[43],c[44],p[23][1],co[234],          s[242],co[237],c[227]);

com4_2 b56(s[57],s[58],s[59],s[60],co[235],             s[243],co[238],c[228]);
com4_2 b57(s[61],s[62],c[45],c[46],co[236],             s[244],co[239],c[229]);
com4_2 b58(c[47],c[48],c[49],c[50],co[237],             s[245],co[240],c[230]);
half_adder b59(p[24][1],p[25][0],                       s[246],co[241]);

com4_2 b60(s[63],s[64],s[65],s[66],co[238],             s[247],co[242],c[231]);
com4_2 b61(s[67],s[68],s[69],c[51],co[239],             s[248],co[243],c[232]);
com4_2 b62(c[52],c[53],c[54],c[55],co[240],             s[249],co[244],c[233]);
full_adder b63(p[26][0],c[56],co[241],                  s[250],co[245]);

com4_2 b64(s[70],s[71],s[72],s[73],co[242],             s[251],co[246],c[234]);
com4_2 b65(s[74],s[75],s[76],c[57],co[243],             s[252],co[247],c[235]);
com4_2 b66(c[58],c[59],c[60],c[61],co[244],             s[253],co[248],c[236]);
full_adder b67(p[27][0],c[62],co[245],                  s[254],co[249]);

com4_2 b68(s[77],s[78],s[79],s[80],co[246],             s[255],co[250],c[237]);
com4_2 b69(s[81],s[82],s[83],c[63],co[247],             s[256],co[251],c[238]);
com4_2 b70(c[64],c[65],c[66],c[67],co[248],             s[257],co[252],c[239]);
com3_2 b71(c[68],c[69],p[28][0],co[249],                s[258],co[253],c[240]);

com4_2 b72(s[84],s[85],s[86],s[87],co[250],            s[259],co[254],c[241]);
com4_2 b73(s[88],s[89],s[90],s[91],co[251],            s[260],co[255],c[242]);
com4_2 b74(c[70],c[71],c[72],c[73],co[252],            s[261],co[256],c[243]);
com3_2 b75(c[74],c[75],c[76],co[253],                  s[262],co[257],c[244]);

com4_2 b76(s[92],s[93],s[94],s[95],co[254],            s[263],co[258],c[245]);
com4_2 b77(s[96],s[97],s[98],s[99],co[255],            s[264],co[259],c[246]);
com4_2 b78(c[77],c[78],c[79],c[80],co[256],            s[265],co[260],c[247]);
com3_2 b79(c[81],c[82],c[83],co[257],            s[266],co[261],c[248]);


com4_2 b80(s[100],s[101],s[102],s[103],co[258],       s[267],co[262],c[249]);
com4_2 b81(s[104],s[105],s[106],s[107],co[259],       s[268],co[263],c[250]);
com4_2 b82(c[85],c[86],c[87],c[88],co[260],           s[269],co[264],c[251]);
com4_2 b83(c[89],c[90],c[91],c[92],co[261],           s[270],co[265],c[252]);

com4_2 b84(s[108],s[109],s[110],s[111],co[262],       s[271],co[266],c[253]);
com4_2 b85(s[112],s[113],s[114],s[115],co[263],       s[272],co[267],c[254]);
com4_2 b86(c[93],c[94],c[95],c[96],co[264],           s[273],co[268],c[255]);
com3_2 b87(c[97],c[98],c[99],co[265],                 s[274],co[269],c[256]);

com4_2 b88(s[116],s[117],s[118],s[119],co[266],       s[275],co[270],c[257]);
com4_2 b89(s[120],s[121],s[122],s[123],co[267],       s[276],co[271],c[258]);
com4_2 b90(c[100],c[101],c[102],c[103],co[268],       s[277],co[272],c[259]);
com3_2 b91(c[104],c[105],c[106],co[269],              s[278],co[273],c[260]);

com4_2 b92(s[124],s[125],s[126],s[127],co[270],       s[279],co[274],c[261]);
com4_2 b93(s[128],s[129],s[130],s[131],co[271],       s[280],co[275],c[262]);
com4_2 b94(c[107],c[108],c[109],c[110],co[272],       s[281],co[276],c[263]);
com3_2 b95(c[111],c[112],c[113],co[273],              s[282],co[277],c[264]);

com4_2 b96(s[132],s[133],s[134],s[135],co[274],       s[283],co[278],c[265]);
com4_2 b97(s[136],s[137],s[138],c[114],co[275],       s[284],co[279],c[266]);
com4_2 b98(c[115],c[116],c[117],c[118],co[276],       s[285],co[280],c[267]);
com4_2 b99(c[119],c[120],c[121],p[31][4],co[277],     s[286],co[281],c[268]);

com4_2 b100(s[139],s[140],s[141],s[142],co[278],      s[287],co[282],c[269]);
com4_2 b101(s[143],s[144],s[145],c[122],co[279],      s[288],co[283],c[270]);
com4_2 b102(c[123],c[124],c[125],c[126],co[280],      s[289],co[284],c[271]);
com3_2 b103(c[127],c[128],p[31][5],co[281],           s[290],co[285],c[272]);

com4_2 b104(s[146],s[147],s[148],s[149],co[282],      s[291],co[286],c[273]);
com4_2 b105(s[150],s[151],c[129],c[130],co[283],      s[292],co[287],c[274]);
com4_2 b106(c[131],c[132],c[133],c[134],co[284],      s[293],co[288],c[275]);
com3_2 b107(c[135],p[31][6],p[30][7],co[285],         s[294],co[289],c[276]);

com4_2 b108(s[152],s[153],s[154],s[155],co[286],      s[295],co[290],c[277]);
com4_2 b109(s[156],s[157],c[136],c[137],co[287],      s[296],co[291],c[278]);
com4_2 b110(c[138],c[139],c[140],c[141],co[288],      s[297],co[292],c[279]);
com3_2 b111(p[31][7],p[30][8],p[29][9],co[289],       s[298],co[293],c[280]);

com4_2 b112(s[158],s[159],s[160],s[161],co[290],      s[299],co[294],c[281]);
com4_2 b113(s[162],c[142],c[143],c[144],co[291],      s[300],co[295],c[282]);
com4_2 b114(c[145],c[146],c[147],p[28][11],co[292],   s[301],co[296],c[283]);
com3_2 b115(p[29][10],p[30][9],p[31][8],co[293],      s[302],co[297],c[284]);

com4_2 b116(s[163],s[164],s[165],s[166],co[294],      s[303],co[298],c[285]);
com4_2 b117(s[167],c[148],c[149],c[150],co[295],      s[304],co[299],c[286]);
com4_2 b118(c[151],c[152],p[27][13],p[28][12],co[296],s[305],co[300],c[287]);
com3_2 b119(p[29][11],p[30][10],p[31][9],co[297],     s[306],co[301],c[288]);

com4_2 b120(s[168],s[169],s[170],s[171],co[298],      s[307],co[302],c[289]);
com4_2 b121(c[153],c[154],c[155],c[156],co[299],      s[308],co[303],c[290]);
com4_2 b122(c[157],p[26][15],p[27][14],p[28][13],co[300],s[309],co[304],c[291]);
com3_2 b123(p[29][12],p[30][11],p[31][10],co[301],      s[310],co[305],c[292]);

com4_2 b124(s[172],s[173],s[174],s[175],co[302],       s[311],co[306],c[293]);
com4_2 b125(c[158],c[159],c[160],c[161],co[303],       s[312],co[307],c[294]);
com4_2 b126(p[25][17],p[26][16],p[27][15],p[28][14],co[304],s[313],co[308],c[295]);
com3_2 b127(p[29][13],p[30][12],p[31][11],co[305],     s[314],co[309],c[296]);

com4_2 b128(s[176],s[178],s[177],c[162],co[306],       s[315],co[310],c[297]);
com4_2 b129(c[163],c[164],c[165],p[24][19],co[307],    s[316],co[311],c[298]);
com4_2 b130(p[25][18],p[26][17],p[27][16],p[28][15],co[308],s[317],co[312],c[299]);
com3_2 b131(p[29][14],p[30][13],p[31][12],co[309],      s[318],co[313],c[300]);

com4_2 b132(s[179],s[180],s[181],c[166],co[310],        s[319],co[314],c[301]);
com4_2 b133(c[167],c[168],p[23][21],p[24][20],co[311],  s[320],co[315],c[302]);
com4_2 b134(p[25][19],p[26][18],p[27][17],p[28][16],co[312],s[321],co[316],c[303]);
com3_2 b135(p[29][15],p[30][14],p[31][13],co[313],      s[322],co[317],c[304]);


com4_2 b136(s[182],s[183],c[169],c[170],co[314],        s[323],co[318],c[305]);
com4_2 b137(c[171],p[22][23],p[23][22],p[24][21],co[315],s[324],co[319],c[306]);
com4_2 b138(p[25][20],p[26][19],p[27][18],p[28][17],co[316],s[325],co[320],c[307]);
com3_2 b139(p[29][16],p[30][15],p[31][14],co[317],         s[326],co[321],c[308]);

com4_2 b140(s[184],s[185],c[172],c[173],co[318],         s[327],co[322],c[309]);
com4_2 b141(p[21][25],p[22][24],p[23][23],p[24][22],co[319],s[328],co[323],c[310]);
com4_2 b142(p[25][21],p[26][20],p[27][19],p[28][18],co[320],s[329],co[324],c[311]);
com3_2 b143(p[29][17],p[30][16],p[31][15],co[321],          s[330],co[325],c[312]);

com4_2 b144(s[186],c[174],c[175],p[20][27],co[322],         s[331],co[326],c[313]);
com4_2 b145(p[21][26],p[22][25],p[23][24],p[24][23],co[323],s[332],co[327],c[314]);
com4_2 b146(p[25][22],p[26][21],p[27][20],p[28][19],co[324],s[333],co[328],c[315]);
com3_2 b147(p[29][18],p[30][17],p[31][16],co[325],          s[334],co[329],c[316]);

com4_2 b148(s[187],c[176],p[19][29],p[20][28],co[326],      s[335],co[330],c[317]);
com4_2 b149(p[21][27],p[22][26],p[23][25],p[24][24],co[327],s[336],co[331],c[318]);
com4_2 b150(p[25][23],p[26][22],p[27][21],p[28][20],co[328],s[337],co[332],c[319]);
com3_2 b151(p[29][19],p[30][18],p[31][17],co[329],          s[338],co[333],c[320]);

com4_2 b152(c[177],p[18][31],p[19][30],p[20][29],co[330],   s[339],co[334],c[321]);
com4_2 b153(p[21][28],p[22][27],p[23][26],p[24][25],co[331],s[340],co[335],c[322]);
com4_2 b154(p[25][24],p[26][23],p[27][22],p[28][21],co[332],s[341],co[336],c[323]);
com3_2 b155(p[29][20],p[30][19],p[31][18],co[333],          s[342],co[337],c[324]);

com4_2 b156(p[19][31],p[20][30],p[21][29],p[22][28],co[334],s[343],co[338],c[325]);
com4_2 b157(p[23][27],p[24][26],p[25][25],p[26][24],co[335],s[344],co[339],c[326]);
com3_2 b158(p[27][23],p[28][22],p[29][21],co[336],          s[345],co[340],c[327]);
full_adder b159(p[30][20],p[31][19],co[337],                s[346],        c[328]);

com4_2 b160(p[20][31],p[21][30],p[22][29],p[23][28],co[338],s[347],co[341],c[329]);
com4_2 b161(p[24][27],p[25][26],p[26][25],p[27][24],co[339],s[348],co[342],c[330]);
com4_2 b162(p[28][23],p[29][22],p[30][21],p[31][20],co[340],s[349],co[343],c[331]);

com4_2 b163(p[21][31],p[22][30],p[23][29],p[24][28],co[341],s[350],co[344],c[332]);
com4_2 b164(p[25][27],p[26][26],p[27][25],p[28][24],co[342],s[351],co[345],c[333]);
com3_2 b165(p[29][23],p[30][22],p[31][21],co[343],          s[352],co[346],c[334]);

com4_2 b166(p[22][31],p[23][30],p[24][29],p[25][28],co[344],s[353],co[347],c[335]);
com4_2 b167(p[26][27],p[27][26],p[28][25],p[29][24],co[345],s[354],co[348],c[336]);
full_adder b168(p[30][23],p[31][22],co[346],                s[355]        ,c[337]);

com4_2 ba167(p[23][31],p[24][30],p[25][29],p[26][28],co[347],s[356],co[349],c[338]);
com3_2 ba168(p[27][27],p[28][26],p[29][25],co[348],          s[357],co[350],c[339]);
half_adder b169(p[30][24],p[31][23],                        s[358],        c[340]);

com4_2 b170(p[24][31],p[25][30],p[26][29],p[27][28],co[349],s[359],co[351],c[341]);
full_adder b171(p[28][27],p[29][26],co[350],                s[360],co[352]);
half_adder b172(p[30][25],p[31][24],                        s[361],        c[342]);

com4_2 b173(p[25][31],p[26][30],p[27][29],p[28][28],co[351],s[362],co[353],c[343]);
com3_2 b174(p[29][27],p[30][26],p[31][25],co[352],          s[363],co[354],c[344]);

com3_2 b175(p[26][31],p[27][30],p[28][29],co[353],          s[364],co[355],c[345]);
com3_2 b176(p[29][28],p[30][27],p[31][26],co[354],          s[365],co[356],c[346]);

com3_2 b177(p[27][31],p[28][30],p[29][29],co[355],          s[366],co[357],c[347]);
full_adder b178(p[30][28],p[31][27],co[356],                s[367],        c[348]);

full_adder b179(p[28][31],p[29][30],co[357],                s[368],        c[349]);
half_adder b180(p[30][29],p[31][28],                        s[369],        c[350]);

half_adder b181(p[29][31],p[30][30],                        s[370],        c[351]);

//stage 3:

assign z[0]=p[0][0];

half_adder c1(p[0][1],p[1][0],          z[1],co[358]);

full_adder c2(s[188],p[2][0],co[358],   z[2],co[359]);

full_adder c3(s[189],p[3][0],co[359],   z[3],co[360]);

com3_2    c4(s[190],c[178],p[4][0],co[360], z[4],co[361],c[352]);

com3_2    c5(s[191],s[192],c[179],co[361],   s[371],co[362],c[353]);

com3_2    c6(s[193],s[194],c[180],co[362],   s[372],co[363],c[354]);

com4_2    c7(s[195],s[196],c[181],c[182],co[363],s[373],co[364],c[355]);

com4_2    c8(s[197],s[198],c[183],c[184],co[364],s[374],co[365],c[356]);

com4_2    c9(s[199],s[200],c[185],c[186],co[365],s[375],co[366],c[357]);

com3_2    c10(s[201],s[202],c[187],co[366],      s[376],co[367],c[358]);
half_adder c11(c[188],p[10][0],                  s[377],co[368]);

com3_2    c12(s[203],s[204],c[189],co[367],      s[378],co[369],c[359]);
full_adder c13(c[190],p[11][0],co[368],          s[379],co[370]);

com3_2    c14(s[205],s[206],c[191],co[369],      s[380],co[371],c[360]);
full_adder c15(c[192],p[12][0],co[370],          s[381],co[372]);

com3_2    c16(s[207],s[208],s[209],co[371],      s[382],co[373],c[361]);
full_adder c17(c[193],c[194],co[372],            s[383],co[374]);

com3_2    c18(s[210],s[211],s[212],co[373],      s[384],co[375],c[362]);
full_adder c19(c[195],c[196],co[374],            s[385],co[376]);

com3_2   c20(s[213],s[214],s[215],co[375],       s[386],co[377],c[363]);
full_adder c21(c[197],c[198],co[376],            s[387],co[378]);

com3_2   c22(s[216],s[217],s[218],co[377],       s[388],co[379],c[364]);
full_adder c23(c[199],c[200],co[378],            s[389],co[380]);

com4_2  c24(s[219],s[220],s[221],c[201],co[379], s[390],co[381],c[365]);
full_adder c25(c[202],c[203],co[380],            s[391],co[382]);

com4_2  c26(s[222],s[223],s[224],c[204],co[381], s[392],co[383],c[366]);
full_adder c27(c[205],c[206],co[382],            s[393],co[384]);

com4_2   c28(s[225],s[226],s[227],c[207],co[383],s[394],co[385],c[367]);
full_adder c29(c[208],c[209],co[384],            s[395],co[386]);

com4_2  c30(s[228],s[229],s[230],c[210],co[385], s[396],co[387],c[368]);
full_adder c31(c[211],c[212],co[386],            s[397],co[388]);

com4_2 c32(s[231],s[232],s[233],c[213],co[387],  s[398],co[389],c[369]);
full_adder c33(c[214],c[215],co[388],            s[399],co[390]);

com4_2  c34(s[234],s[235],s[236],c[216],co[389], s[400],co[391],c[370]);
com3_2  c35(c[217],c[218],p[22][0],co[390],      s[401],co[392],c[371]);

com4_2  c36(s[237],s[238],s[239],c[219],co[391], s[402],co[393],c[372]);
com3_2  c37(c[220],c[221],p[23][0],co[392],      s[403],co[394],c[373]);

com4_2 c38(s[240],s[241],s[242],c[222],co[393],  s[404],co[395],c[374]);
com3_2 c39(c[223],c[224],p[24][0],co[394],       s[405],co[396],c[375]);

com4_2 c40(s[243],s[244],s[245],s[246],co[395],  s[406],co[397],c[376]);
com3_2 c41(c[225],c[226],c[227],co[396],         s[407],co[398],c[377]);

com4_2 c42(s[247],s[248],s[249],s[250],co[397],  s[408],co[399],c[378]);
com3_2 c43(c[228],c[229],c[230],co[398],         s[409],co[400],c[379]);

com4_2 c44(s[251],s[252],s[253],s[254],co[399],  s[410],co[401],c[380]);
com3_2 c45(c[231],c[232],c[233],co[400],         s[411],co[402],c[381]);

com4_2 c46(s[255],s[256],s[257],s[258],co[401],  s[412],co[403],c[382]);
com3_2 c47(c[234],c[235],c[236],co[402],         s[413],co[404],c[383]);

com4_2 c48(s[259],s[260],s[261],s[262],co[403],  s[414],co[405],c[384]);
com4_2 c49(c[237],c[238],c[239],c[240],co[404],  s[415],co[406],c[385]);

com4_2 c50(s[263],s[264],s[265],s[266],co[405],  s[416],co[407],c[386]);
com4_2 c51(c[241],c[242],c[243],c[244],co[406],  s[417],co[408],c[387]);

com4_2 c52(s[267],s[268],s[269],s[270],co[407],  s[418],co[409],c[388]);
com4_2 c53(c[245],c[246],c[247],c[248],co[408],  s[419],co[410],c[389]);

com4_2 c54(s[271],s[272],s[273],s[274],co[409],  s[420],co[411],c[390]);
com4_2 c55(c[249],c[250],c[251],c[252],co[410],  s[421],co[412],c[391]);

com4_2 c56(s[275],s[276],s[277],s[278],co[411],  s[422],co[413],c[392]);
com4_2 c57(c[253],c[254],c[255],c[256],co[412],  s[423],co[414],c[393]);

com4_2 c58(s[279],s[280],s[281],s[282],co[413],  s[424],co[415],c[394]);
com4_2 c59(c[257],c[258],c[259],c[260],co[414],  s[425],co[416],c[395]);

com4_2 c60(s[283],s[284],s[285],s[286],co[415],  s[426],co[417],c[396]);
com4_2 c61(c[261],c[262],c[263],c[264],co[416],  s[427],co[418],c[397]);

com4_2 c62(s[287],s[288],s[289],s[290],co[417],  s[428],co[419],c[398]);
com4_2 c63(c[265],c[266],c[267],c[268],co[418],  s[429],co[420],c[399]);

com4_2 c64(s[291],s[292],s[293],s[294],co[419],  s[430],co[421],c[400]);
com4_2 c65(c[269],c[270],c[271],c[272],co[420],  s[431],co[422],c[401]);

com4_2 c66(s[295],s[296],s[297],s[298],co[421],  s[432],co[423],c[402]);
com4_2 c67(c[273],c[274],c[275],c[276],co[422],  s[433],co[424],c[403]);

com4_2 c68(s[299],s[300],s[301],s[302],co[423],  s[434],co[425],c[404]);
com4_2 c69(c[277],c[278],c[279],c[280],co[424],  s[435],co[426],c[405]);

com4_2 c70(s[303],s[304],s[305],s[306],co[425],  s[436],co[427],c[406]);
com4_2 c71(c[281],c[282],c[283],c[284],co[426],  s[437],co[428],c[407]);

com4_2 c72(s[307],s[308],s[309],s[310],co[427],  s[438],co[429],c[408]);
com4_2 c73(c[285],c[286],c[287],c[288],co[428],  s[439],co[430],c[409]);

com4_2 c74(s[311],s[312],s[313],s[314],co[429],  s[440],co[431],c[410]);
com4_2 c75(c[289],c[290],c[291],c[292],co[430],  s[441],co[432],c[411]);

com4_2 c76(s[315],s[316],s[317],s[318],co[431],  s[442],co[433],c[412]);
com4_2 c77(c[293],c[294],c[295],c[296],co[432],  s[443],co[434],c[413]);

com4_2 c78(s[319],s[320],s[321],s[322],co[433],  s[444],co[435],c[414]);
com4_2 c79(c[297],c[298],c[299],c[300],co[434],  s[445],co[436],c[415]);

com4_2 c80(s[323],s[324],s[325],s[326],co[435],  s[446],co[437],c[416]);
com4_2 c81(c[301],c[302],c[303],c[304],co[436],  s[447],co[438],c[417]);

com4_2 c82(s[327],s[328],s[329],s[330],co[437],  s[448],co[439],c[418]);
com4_2 c83(c[305],c[306],c[307],c[308],co[438],  s[449],co[440],c[419]);

com4_2 c84(s[331],s[332],s[333],s[334],co[439],  s[450],co[441],c[420]);
com4_2 c85(c[309],c[310],c[311],c[312],co[440],  s[451],co[442],c[421]);

com4_2 c86(s[335],s[336],s[337],s[338],co[441],  s[452],co[443],c[422]);
com4_2 c87(c[313],c[314],c[315],c[316],co[442],  s[453],co[444],c[423]);

com4_2 c88(s[339],s[340],s[341],s[342],co[443],  s[454],co[445],c[424]);
com4_2 c89(c[317],c[318],c[319],c[320],co[444],  s[455],co[446],c[425]);

com4_2 c90(s[343],s[344],s[345],s[346],co[445],  s[456],co[447],c[426]);
com4_2 c91(c[321],c[322],c[323],c[324],co[446],  s[457],co[448],c[427]);

com4_2 c92(s[347],s[348],s[349],c[325],co[447],  s[458],co[449],c[428]);
com3_2 c93(c[326],c[327],c[328],co[448],         s[459],co[450],c[429]);

com4_2 c94(s[350],s[351],s[352],c[329],co[449],  s[460],co[451],c[430]);
full_adder c95(c[330],c[331],co[450],            s[461],co[452]);

com4_2 c96(s[353],s[354],s[355],c[332],co[451],  s[462],co[453],c[431]);
full_adder c97(c[333],c[334],co[452],            s[463],co[454]);

com4_2 c98(s[356],s[357],s[358],c[335],co[453],  s[464],co[455],c[432]);
full_adder c99(c[336],c[337],co[454],            s[465],co[456]);

com4_2 d1(s[359],s[360],s[361],c[338],co[455],   s[466],co[457],c[433]);
full_adder d2(c[339],c[340],co[456],             s[467],co[458]);

full_adder d3(s[362],s[363],co[457],             s[468],co[459]);
full_adder d4(c[341],c[342],co[458],             s[469],co[460]);

full_adder d5(s[364],s[365],co[459],             s[470],co[461]);
full_adder d6(c[343],c[344],co[460],             s[471],co[462]);

full_adder d7(s[366],s[367],co[461],             s[472],co[463]);
full_adder d8(c[345],c[346],co[462],             s[473],co[464]);

full_adder d9(s[368],s[369],co[463],             s[474],co[465]);
full_adder d10(c[347],c[348],co[464],            s[475],co[466]);

full_adder d11(s[370],c[349],co[465],            s[476],co[467]);
full_adder d12(c[350],p[31][29],co[466],         s[477],co[468]);

full_adder d13(c[351],p[30][31],co[467],         s[478],co[469]);
half_adder d14(p[31][30],co[468],                s[479],co[470]);

full_adder d15(p[31][31],co[469],co[470],        s[480],c[435]);

//stage 4:

half_adder q1(c[352],s[371],                      z[5],  co[471]);
full_adder q2(c[353],s[372],              co[471],z[6],  co[472]);
full_adder q3(c[354],s[373],              co[472],z[7],  co[473]);
full_adder q4(c[355],s[374],              co[473],z[8],  co[474]);
full_adder q5(c[356],s[375],              co[474],z[9],  co[475]);
com3_2     q6(c[357],s[376],s[377],       co[475],z[10], co[476],c[436]);
com3_2     q7(c[358],s[378],s[379],       co[476],s[481],co[477],c[437]);
com3_2     q8(c[359],s[380],s[381],       co[477],s[482],co[478],c[438]);
com3_2     q9(c[360],s[382],s[383],       co[478],s[483],co[479],c[439]);
com3_2    q10(c[361],s[384],s[385],       co[479],s[484],co[480],c[440]);
com3_2    q11(c[362],s[386],s[387],       co[480],s[485],co[481],c[441]);
com3_2    q12(c[363],s[388],s[389],       co[481],s[486],co[482],c[442]);
com3_2    q13(c[364],s[390],s[391],       co[482],s[487],co[483],c[443]);
com3_2    q14(c[365],s[392],s[393],       co[483],s[488],co[484],c[444]);
com3_2    q15(c[366],s[394],s[395],       co[484],s[489],co[485],c[445]);
com3_2    q16(c[367],s[396],s[397],       co[485],s[490],co[486],c[446]);
com3_2    q17(c[368],s[398],s[399],       co[486],s[491],co[487],c[447]);
com3_2    q18(c[369],s[400],s[401],       co[487],s[492],co[488],c[448]);
com4_2    q19(c[370],c[371],s[402],s[403],co[488],s[493],co[489],c[449]);
com4_2    q20(c[372],c[373],s[404],s[405],co[489],s[494],co[490],c[450]);
com4_2    q21(c[374],c[375],s[406],s[407],co[490],s[495],co[491],c[451]);
com4_2    q22(c[376],c[377],s[408],s[409],co[491],s[496],co[492],c[452]);
com4_2    q23(c[378],c[379],s[410],s[411],co[492],s[497],co[493],c[453]);
com4_2    q24(c[380],c[381],s[412],s[413],co[493],s[498],co[494],c[454]);
com4_2    q25(c[382],c[383],s[414],s[415],co[494],s[499],co[495],c[455]);
com4_2    q26(c[384],c[385],s[416],s[417],co[495],s[500],co[496],c[456]);
com4_2    q27(c[386],c[387],s[418],s[419],co[496],s[501],co[497],c[457]);
com4_2    q28(c[388],c[389],s[420],s[421],co[497],s[502],co[498],c[458]);
com4_2    q29(c[390],c[391],s[422],s[423],co[498],s[503],co[499],c[459]);
com4_2    q30(c[392],c[393],s[424],s[425],co[499],s[504],co[500],c[460]);
com4_2    q31(c[394],c[395],s[426],s[427],co[500],s[505],co[501],c[461]);
com4_2    q32(c[396],c[397],s[428],s[429],co[501],s[506],co[502],c[462]);
com4_2    q33(c[398],c[399],s[430],s[431],co[502],s[507],co[503],c[463]);
com4_2    q34(c[400],c[401],s[432],s[433],co[503],s[508],co[504],c[464]);
com4_2    q35(c[402],c[403],s[434],s[435],co[504],s[509],co[505],c[465]);
com4_2    q36(c[404],c[405],s[436],s[437],co[505],s[510],co[506],c[466]);
com4_2    q37(c[406],c[407],s[438],s[439],co[506],s[511],co[507],c[467]);
com4_2    q38(c[408],c[409],s[440],s[441],co[507],s[512],co[508],c[468]);
com4_2    q39(c[410],c[411],s[442],s[443],co[508],s[513],co[509],c[469]);
com4_2    q40(c[412],c[413],s[444],s[445],co[509],s[514],co[510],c[470]);
com4_2    q41(c[414],c[415],s[446],s[447],co[510],s[515],co[511],c[471]);
com4_2    q42(c[416],c[417],s[448],s[449],co[511],s[516],co[512],c[472]);
com4_2    q43(c[418],c[419],s[450],s[451],co[512],s[517],co[513],c[473]);
com4_2    q44(c[420],c[421],s[452],s[453],co[513],s[518],co[514],c[474]);
com4_2    q45(c[422],c[423],s[454],s[455],co[514],s[519],co[515],c[475]);
com4_2    q46(c[424],c[425],s[456],s[457],co[515],s[520],co[516],c[476]);
com4_2    q47(c[426],c[427],s[458],s[459],co[516],s[521],co[517],c[477]);
com4_2    q48(c[428],c[429],s[460],s[461],co[517],s[522],co[518],c[478]);
com3_2    q49(c[430],s[462],s[463],       co[518],s[523],co[519],c[479]);
com3_2    q50(c[431],s[464],s[465],       co[519],s[524],co[520],c[480]);
com3_2    q51(c[432],s[466],s[467],       co[520],s[525],co[521],c[481]);
com3_2    q52(c[433],s[468],s[469],       co[521],s[526],co[522],c[482]);
full_adder q53(      s[470],s[471],       co[522],s[527],co[523]);
full_adder q54(      s[472],s[473],       co[523],s[528],co[524]);
full_adder q55(      s[474],s[475],       co[524],s[529],co[525]);
full_adder q56(      s[476],s[477],       co[525],s[530],co[526]);
full_adder q57(      s[478],s[479],       co[526],s[531],        c[483]);


half_adder w1( c[436],s[481],        z[11],co[527]);
full_adder w2( c[437],s[482],co[527],z[12],co[528]);
full_adder w3( c[438],s[483],co[528],z[13],co[529]);
full_adder w4( c[439],s[484],co[529],z[14],co[530]);
full_adder w5( c[440],s[485],co[530],z[15],co[531]);
full_adder w6( c[441],s[486],co[531],z[16],co[532]);
full_adder w7( c[442],s[487],co[532],z[17],co[533]);
full_adder w8( c[443],s[488],co[533],z[18],co[534]);
full_adder w9( c[444],s[489],co[534],z[19],co[535]);
full_adder w10(c[445],s[490],co[535],z[20],co[536]);
full_adder w11(c[446],s[491],co[536],z[21],co[537]);
full_adder w12(c[447],s[492],co[537],z[22],co[538]);
full_adder w13(c[448],s[493],co[538],z[23],co[539]);
full_adder w14(c[449],s[494],co[539],z[24],co[540]);
full_adder w15(c[450],s[495],co[540],z[25],co[541]);
full_adder w16(c[451],s[496],co[541],z[26],co[542]);
full_adder w17(c[452],s[497],co[542],z[27],co[543]);
full_adder w18(c[453],s[498],co[543],z[28],co[544]);
full_adder w19(c[454],s[499],co[544],z[29],co[545]);
full_adder w20(c[455],s[500],co[545],z[30],co[546]);
full_adder w21(c[456],s[501],co[546],z[31],co[547]);
full_adder w22(c[457],s[502],co[547],z[32],co[548]);
full_adder w23(c[458],s[503],co[548],z[33],co[549]);
full_adder w24(c[459],s[504],co[549],z[34],co[550]);
full_adder w25(c[460],s[505],co[550],z[35],co[551]);
full_adder w26(c[461],s[506],co[551],z[36],co[552]);
full_adder w27(c[462],s[507],co[552],z[37],co[553]);
full_adder w28(c[463],s[508],co[553],z[38],co[554]);
full_adder w29(c[464],s[509],co[554],z[39],co[555]);
full_adder w30(c[465],s[510],co[555],z[40],co[556]);
full_adder w31(c[466],s[511],co[556],z[41],co[557]);
full_adder w32(c[467],s[512],co[557],z[42],co[558]);
full_adder w33(c[468],s[513],co[558],z[43],co[559]);
full_adder w34(c[469],s[514],co[559],z[44],co[560]);
full_adder w35(c[470],s[515],co[560],z[45],co[561]);
full_adder w36(c[471],s[516],co[561],z[46],co[562]);
full_adder w37(c[472],s[517],co[562],z[47],co[563]);
full_adder w38(c[473],s[518],co[563],z[48],co[564]);
full_adder w39(c[474],s[519],co[564],z[49],co[565]);
full_adder w40(c[475],s[520],co[565],z[50],co[566]);
full_adder w41(c[476],s[521],co[566],z[51],co[567]);
full_adder w42(c[477],s[522],co[567],z[52],co[568]);
full_adder w43(c[478],s[523],co[568],z[53],co[569]);
full_adder w44(c[479],s[524],co[569],z[54],co[570]);
full_adder w45(c[480],s[525],co[570],z[55],co[571]);
full_adder w46(c[481],s[526],co[571],z[56],co[572]);
full_adder w47(c[482],s[527],co[572],z[57],co[573]);
half_adder w48(       s[528],co[573],z[58],co[574]);
half_adder w49(       s[529],co[574],z[59],co[575]);
half_adder w50(       s[530],co[575],z[60],co[576]);
half_adder w51(       s[531],co[576],z[61],co[577]);
full_adder w52(c[483],s[480],co[577],z[62],co[578]);
half_adder w53(c[435],       co[578],z[63],co[579]);







endmodule
